** Profile: "Plan A DC-DC Test"  [ F:\Programs\Verilog\FPGA_Group\test_br0101\analog\br0101_ad9239\br0101_ad9239-pspicefiles\plan a dc\dc test.sim ] 

** Creating circuit file "DC Test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "F:/Programs/Verilog/FPGA_Group/test_br0101/analog/br0101_ad9286/models/ada4937.lib" 
* From [PSPICE NETLIST] section of G:\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.0.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_Vi -3.63 3.67 0.05 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Plan A DC.net" 


.END
