//-----------------------------------------------------------------------------
// lmb_bram_elaborate.v
//-----------------------------------------------------------------------------

`timescale 1 ps / 100 fs

`uselib lib=unisims_ver

module lmb_bram_elaborate
  (
    BRAM_Rst_A,
    BRAM_Clk_A,
    BRAM_EN_A,
    BRAM_WEN_A,
    BRAM_Addr_A,
    BRAM_Din_A,
    BRAM_Dout_A,
    BRAM_Rst_B,
    BRAM_Clk_B,
    BRAM_EN_B,
    BRAM_WEN_B,
    BRAM_Addr_B,
    BRAM_Din_B,
    BRAM_Dout_B
  );
  parameter
    C_MEMSIZE = 'h10000,
    C_PORT_DWIDTH = 32,
    C_PORT_AWIDTH = 32,
    C_NUM_WE = 4,
    C_FAMILY = "virtex4";
  input BRAM_Rst_A;
  input BRAM_Clk_A;
  input BRAM_EN_A;
  input [0:C_NUM_WE-1] BRAM_WEN_A;
  input [0:C_PORT_AWIDTH-1] BRAM_Addr_A;
  output [0:C_PORT_DWIDTH-1] BRAM_Din_A;
  input [0:C_PORT_DWIDTH-1] BRAM_Dout_A;
  input BRAM_Rst_B;
  input BRAM_Clk_B;
  input BRAM_EN_B;
  input [0:C_NUM_WE-1] BRAM_WEN_B;
  input [0:C_PORT_AWIDTH-1] BRAM_Addr_B;
  output [0:C_PORT_DWIDTH-1] BRAM_Din_B;
  input [0:C_PORT_DWIDTH-1] BRAM_Dout_B;

  // Internal signals

  wire net_gnd0;
  wire [3:0] net_gnd4;
  wire [0:0] pgassign1;
  wire [0:30] pgassign2;
  wire [14:0] pgassign3;
  wire [31:0] pgassign4;
  wire [31:0] pgassign5;
  wire [3:0] pgassign6;
  wire [14:0] pgassign7;
  wire [31:0] pgassign8;
  wire [31:0] pgassign9;
  wire [3:0] pgassign10;
  wire [14:0] pgassign11;
  wire [31:0] pgassign12;
  wire [31:0] pgassign13;
  wire [3:0] pgassign14;
  wire [14:0] pgassign15;
  wire [31:0] pgassign16;
  wire [31:0] pgassign17;
  wire [3:0] pgassign18;
  wire [14:0] pgassign19;
  wire [31:0] pgassign20;
  wire [31:0] pgassign21;
  wire [3:0] pgassign22;
  wire [14:0] pgassign23;
  wire [31:0] pgassign24;
  wire [31:0] pgassign25;
  wire [3:0] pgassign26;
  wire [14:0] pgassign27;
  wire [31:0] pgassign28;
  wire [31:0] pgassign29;
  wire [3:0] pgassign30;
  wire [14:0] pgassign31;
  wire [31:0] pgassign32;
  wire [31:0] pgassign33;
  wire [3:0] pgassign34;
  wire [14:0] pgassign35;
  wire [31:0] pgassign36;
  wire [31:0] pgassign37;
  wire [3:0] pgassign38;
  wire [14:0] pgassign39;
  wire [31:0] pgassign40;
  wire [31:0] pgassign41;
  wire [3:0] pgassign42;
  wire [14:0] pgassign43;
  wire [31:0] pgassign44;
  wire [31:0] pgassign45;
  wire [3:0] pgassign46;
  wire [14:0] pgassign47;
  wire [31:0] pgassign48;
  wire [31:0] pgassign49;
  wire [3:0] pgassign50;
  wire [14:0] pgassign51;
  wire [31:0] pgassign52;
  wire [31:0] pgassign53;
  wire [3:0] pgassign54;
  wire [14:0] pgassign55;
  wire [31:0] pgassign56;
  wire [31:0] pgassign57;
  wire [3:0] pgassign58;
  wire [14:0] pgassign59;
  wire [31:0] pgassign60;
  wire [31:0] pgassign61;
  wire [3:0] pgassign62;
  wire [14:0] pgassign63;
  wire [31:0] pgassign64;
  wire [31:0] pgassign65;
  wire [3:0] pgassign66;
  wire [14:0] pgassign67;
  wire [31:0] pgassign68;
  wire [31:0] pgassign69;
  wire [3:0] pgassign70;
  wire [14:0] pgassign71;
  wire [31:0] pgassign72;
  wire [31:0] pgassign73;
  wire [3:0] pgassign74;
  wire [14:0] pgassign75;
  wire [31:0] pgassign76;
  wire [31:0] pgassign77;
  wire [3:0] pgassign78;
  wire [14:0] pgassign79;
  wire [31:0] pgassign80;
  wire [31:0] pgassign81;
  wire [3:0] pgassign82;
  wire [14:0] pgassign83;
  wire [31:0] pgassign84;
  wire [31:0] pgassign85;
  wire [3:0] pgassign86;
  wire [14:0] pgassign87;
  wire [31:0] pgassign88;
  wire [31:0] pgassign89;
  wire [3:0] pgassign90;
  wire [14:0] pgassign91;
  wire [31:0] pgassign92;
  wire [31:0] pgassign93;
  wire [3:0] pgassign94;
  wire [14:0] pgassign95;
  wire [31:0] pgassign96;
  wire [31:0] pgassign97;
  wire [3:0] pgassign98;
  wire [14:0] pgassign99;
  wire [31:0] pgassign100;
  wire [31:0] pgassign101;
  wire [3:0] pgassign102;
  wire [14:0] pgassign103;
  wire [31:0] pgassign104;
  wire [31:0] pgassign105;
  wire [3:0] pgassign106;
  wire [14:0] pgassign107;
  wire [31:0] pgassign108;
  wire [31:0] pgassign109;
  wire [3:0] pgassign110;
  wire [14:0] pgassign111;
  wire [31:0] pgassign112;
  wire [31:0] pgassign113;
  wire [3:0] pgassign114;
  wire [14:0] pgassign115;
  wire [31:0] pgassign116;
  wire [31:0] pgassign117;
  wire [3:0] pgassign118;
  wire [14:0] pgassign119;
  wire [31:0] pgassign120;
  wire [31:0] pgassign121;
  wire [3:0] pgassign122;
  wire [14:0] pgassign123;
  wire [31:0] pgassign124;
  wire [31:0] pgassign125;
  wire [3:0] pgassign126;
  wire [14:0] pgassign127;
  wire [31:0] pgassign128;
  wire [31:0] pgassign129;
  wire [3:0] pgassign130;
  wire [14:0] pgassign131;
  wire [31:0] pgassign132;
  wire [31:0] pgassign133;
  wire [3:0] pgassign134;
  wire [14:0] pgassign135;
  wire [31:0] pgassign136;
  wire [31:0] pgassign137;
  wire [3:0] pgassign138;
  wire [14:0] pgassign139;
  wire [31:0] pgassign140;
  wire [31:0] pgassign141;
  wire [3:0] pgassign142;
  wire [14:0] pgassign143;
  wire [31:0] pgassign144;
  wire [31:0] pgassign145;
  wire [3:0] pgassign146;
  wire [14:0] pgassign147;
  wire [31:0] pgassign148;
  wire [31:0] pgassign149;
  wire [3:0] pgassign150;
  wire [14:0] pgassign151;
  wire [31:0] pgassign152;
  wire [31:0] pgassign153;
  wire [3:0] pgassign154;
  wire [14:0] pgassign155;
  wire [31:0] pgassign156;
  wire [31:0] pgassign157;
  wire [3:0] pgassign158;
  wire [14:0] pgassign159;
  wire [31:0] pgassign160;
  wire [31:0] pgassign161;
  wire [3:0] pgassign162;
  wire [14:0] pgassign163;
  wire [31:0] pgassign164;
  wire [31:0] pgassign165;
  wire [3:0] pgassign166;
  wire [14:0] pgassign167;
  wire [31:0] pgassign168;
  wire [31:0] pgassign169;
  wire [3:0] pgassign170;
  wire [14:0] pgassign171;
  wire [31:0] pgassign172;
  wire [31:0] pgassign173;
  wire [3:0] pgassign174;
  wire [14:0] pgassign175;
  wire [31:0] pgassign176;
  wire [31:0] pgassign177;
  wire [3:0] pgassign178;
  wire [14:0] pgassign179;
  wire [31:0] pgassign180;
  wire [31:0] pgassign181;
  wire [3:0] pgassign182;
  wire [14:0] pgassign183;
  wire [31:0] pgassign184;
  wire [31:0] pgassign185;
  wire [3:0] pgassign186;
  wire [14:0] pgassign187;
  wire [31:0] pgassign188;
  wire [31:0] pgassign189;
  wire [3:0] pgassign190;
  wire [14:0] pgassign191;
  wire [31:0] pgassign192;
  wire [31:0] pgassign193;
  wire [3:0] pgassign194;
  wire [14:0] pgassign195;
  wire [31:0] pgassign196;
  wire [31:0] pgassign197;
  wire [3:0] pgassign198;
  wire [14:0] pgassign199;
  wire [31:0] pgassign200;
  wire [31:0] pgassign201;
  wire [3:0] pgassign202;
  wire [14:0] pgassign203;
  wire [31:0] pgassign204;
  wire [31:0] pgassign205;
  wire [3:0] pgassign206;
  wire [14:0] pgassign207;
  wire [31:0] pgassign208;
  wire [31:0] pgassign209;
  wire [3:0] pgassign210;
  wire [14:0] pgassign211;
  wire [31:0] pgassign212;
  wire [31:0] pgassign213;
  wire [3:0] pgassign214;
  wire [14:0] pgassign215;
  wire [31:0] pgassign216;
  wire [31:0] pgassign217;
  wire [3:0] pgassign218;
  wire [14:0] pgassign219;
  wire [31:0] pgassign220;
  wire [31:0] pgassign221;
  wire [3:0] pgassign222;
  wire [14:0] pgassign223;
  wire [31:0] pgassign224;
  wire [31:0] pgassign225;
  wire [3:0] pgassign226;
  wire [14:0] pgassign227;
  wire [31:0] pgassign228;
  wire [31:0] pgassign229;
  wire [3:0] pgassign230;
  wire [14:0] pgassign231;
  wire [31:0] pgassign232;
  wire [31:0] pgassign233;
  wire [3:0] pgassign234;
  wire [14:0] pgassign235;
  wire [31:0] pgassign236;
  wire [31:0] pgassign237;
  wire [3:0] pgassign238;
  wire [14:0] pgassign239;
  wire [31:0] pgassign240;
  wire [31:0] pgassign241;
  wire [3:0] pgassign242;
  wire [14:0] pgassign243;
  wire [31:0] pgassign244;
  wire [31:0] pgassign245;
  wire [3:0] pgassign246;
  wire [14:0] pgassign247;
  wire [31:0] pgassign248;
  wire [31:0] pgassign249;
  wire [3:0] pgassign250;
  wire [14:0] pgassign251;
  wire [31:0] pgassign252;
  wire [31:0] pgassign253;
  wire [3:0] pgassign254;
  wire [14:0] pgassign255;
  wire [31:0] pgassign256;
  wire [31:0] pgassign257;
  wire [3:0] pgassign258;

  // Internal assignments

  assign pgassign1[0:0] = 1'b1;
  assign pgassign2[0:30] = 31'b0000000000000000000000000000000;
  assign pgassign3[14:14] = 1'b1;
  assign pgassign3[13:0] = BRAM_Addr_A[16:29];
  assign pgassign4[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign4[0:0] = BRAM_Dout_A[0:0];
  assign BRAM_Din_A[0:0] = pgassign5[0:0];
  assign pgassign6[3:3] = BRAM_WEN_A[0:0];
  assign pgassign6[2:2] = BRAM_WEN_A[0:0];
  assign pgassign6[1:1] = BRAM_WEN_A[0:0];
  assign pgassign6[0:0] = BRAM_WEN_A[0:0];
  assign pgassign7[14:14] = 1'b1;
  assign pgassign7[13:0] = BRAM_Addr_B[16:29];
  assign pgassign8[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign8[0:0] = BRAM_Dout_B[0:0];
  assign BRAM_Din_B[0:0] = pgassign9[0:0];
  assign pgassign10[3:3] = BRAM_WEN_B[0:0];
  assign pgassign10[2:2] = BRAM_WEN_B[0:0];
  assign pgassign10[1:1] = BRAM_WEN_B[0:0];
  assign pgassign10[0:0] = BRAM_WEN_B[0:0];
  assign pgassign11[14:14] = 1'b1;
  assign pgassign11[13:0] = BRAM_Addr_A[16:29];
  assign pgassign12[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign12[0:0] = BRAM_Dout_A[1:1];
  assign BRAM_Din_A[1:1] = pgassign13[0:0];
  assign pgassign14[3:3] = BRAM_WEN_A[0:0];
  assign pgassign14[2:2] = BRAM_WEN_A[0:0];
  assign pgassign14[1:1] = BRAM_WEN_A[0:0];
  assign pgassign14[0:0] = BRAM_WEN_A[0:0];
  assign pgassign15[14:14] = 1'b1;
  assign pgassign15[13:0] = BRAM_Addr_B[16:29];
  assign pgassign16[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign16[0:0] = BRAM_Dout_B[1:1];
  assign BRAM_Din_B[1:1] = pgassign17[0:0];
  assign pgassign18[3:3] = BRAM_WEN_B[0:0];
  assign pgassign18[2:2] = BRAM_WEN_B[0:0];
  assign pgassign18[1:1] = BRAM_WEN_B[0:0];
  assign pgassign18[0:0] = BRAM_WEN_B[0:0];
  assign pgassign19[14:14] = 1'b1;
  assign pgassign19[13:0] = BRAM_Addr_A[16:29];
  assign pgassign20[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign20[0:0] = BRAM_Dout_A[2:2];
  assign BRAM_Din_A[2:2] = pgassign21[0:0];
  assign pgassign22[3:3] = BRAM_WEN_A[0:0];
  assign pgassign22[2:2] = BRAM_WEN_A[0:0];
  assign pgassign22[1:1] = BRAM_WEN_A[0:0];
  assign pgassign22[0:0] = BRAM_WEN_A[0:0];
  assign pgassign23[14:14] = 1'b1;
  assign pgassign23[13:0] = BRAM_Addr_B[16:29];
  assign pgassign24[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign24[0:0] = BRAM_Dout_B[2:2];
  assign BRAM_Din_B[2:2] = pgassign25[0:0];
  assign pgassign26[3:3] = BRAM_WEN_B[0:0];
  assign pgassign26[2:2] = BRAM_WEN_B[0:0];
  assign pgassign26[1:1] = BRAM_WEN_B[0:0];
  assign pgassign26[0:0] = BRAM_WEN_B[0:0];
  assign pgassign27[14:14] = 1'b1;
  assign pgassign27[13:0] = BRAM_Addr_A[16:29];
  assign pgassign28[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign28[0:0] = BRAM_Dout_A[3:3];
  assign BRAM_Din_A[3:3] = pgassign29[0:0];
  assign pgassign30[3:3] = BRAM_WEN_A[0:0];
  assign pgassign30[2:2] = BRAM_WEN_A[0:0];
  assign pgassign30[1:1] = BRAM_WEN_A[0:0];
  assign pgassign30[0:0] = BRAM_WEN_A[0:0];
  assign pgassign31[14:14] = 1'b1;
  assign pgassign31[13:0] = BRAM_Addr_B[16:29];
  assign pgassign32[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign32[0:0] = BRAM_Dout_B[3:3];
  assign BRAM_Din_B[3:3] = pgassign33[0:0];
  assign pgassign34[3:3] = BRAM_WEN_B[0:0];
  assign pgassign34[2:2] = BRAM_WEN_B[0:0];
  assign pgassign34[1:1] = BRAM_WEN_B[0:0];
  assign pgassign34[0:0] = BRAM_WEN_B[0:0];
  assign pgassign35[14:14] = 1'b1;
  assign pgassign35[13:0] = BRAM_Addr_A[16:29];
  assign pgassign36[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign36[0:0] = BRAM_Dout_A[4:4];
  assign BRAM_Din_A[4:4] = pgassign37[0:0];
  assign pgassign38[3:3] = BRAM_WEN_A[0:0];
  assign pgassign38[2:2] = BRAM_WEN_A[0:0];
  assign pgassign38[1:1] = BRAM_WEN_A[0:0];
  assign pgassign38[0:0] = BRAM_WEN_A[0:0];
  assign pgassign39[14:14] = 1'b1;
  assign pgassign39[13:0] = BRAM_Addr_B[16:29];
  assign pgassign40[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign40[0:0] = BRAM_Dout_B[4:4];
  assign BRAM_Din_B[4:4] = pgassign41[0:0];
  assign pgassign42[3:3] = BRAM_WEN_B[0:0];
  assign pgassign42[2:2] = BRAM_WEN_B[0:0];
  assign pgassign42[1:1] = BRAM_WEN_B[0:0];
  assign pgassign42[0:0] = BRAM_WEN_B[0:0];
  assign pgassign43[14:14] = 1'b1;
  assign pgassign43[13:0] = BRAM_Addr_A[16:29];
  assign pgassign44[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign44[0:0] = BRAM_Dout_A[5:5];
  assign BRAM_Din_A[5:5] = pgassign45[0:0];
  assign pgassign46[3:3] = BRAM_WEN_A[0:0];
  assign pgassign46[2:2] = BRAM_WEN_A[0:0];
  assign pgassign46[1:1] = BRAM_WEN_A[0:0];
  assign pgassign46[0:0] = BRAM_WEN_A[0:0];
  assign pgassign47[14:14] = 1'b1;
  assign pgassign47[13:0] = BRAM_Addr_B[16:29];
  assign pgassign48[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign48[0:0] = BRAM_Dout_B[5:5];
  assign BRAM_Din_B[5:5] = pgassign49[0:0];
  assign pgassign50[3:3] = BRAM_WEN_B[0:0];
  assign pgassign50[2:2] = BRAM_WEN_B[0:0];
  assign pgassign50[1:1] = BRAM_WEN_B[0:0];
  assign pgassign50[0:0] = BRAM_WEN_B[0:0];
  assign pgassign51[14:14] = 1'b1;
  assign pgassign51[13:0] = BRAM_Addr_A[16:29];
  assign pgassign52[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign52[0:0] = BRAM_Dout_A[6:6];
  assign BRAM_Din_A[6:6] = pgassign53[0:0];
  assign pgassign54[3:3] = BRAM_WEN_A[0:0];
  assign pgassign54[2:2] = BRAM_WEN_A[0:0];
  assign pgassign54[1:1] = BRAM_WEN_A[0:0];
  assign pgassign54[0:0] = BRAM_WEN_A[0:0];
  assign pgassign55[14:14] = 1'b1;
  assign pgassign55[13:0] = BRAM_Addr_B[16:29];
  assign pgassign56[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign56[0:0] = BRAM_Dout_B[6:6];
  assign BRAM_Din_B[6:6] = pgassign57[0:0];
  assign pgassign58[3:3] = BRAM_WEN_B[0:0];
  assign pgassign58[2:2] = BRAM_WEN_B[0:0];
  assign pgassign58[1:1] = BRAM_WEN_B[0:0];
  assign pgassign58[0:0] = BRAM_WEN_B[0:0];
  assign pgassign59[14:14] = 1'b1;
  assign pgassign59[13:0] = BRAM_Addr_A[16:29];
  assign pgassign60[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign60[0:0] = BRAM_Dout_A[7:7];
  assign BRAM_Din_A[7:7] = pgassign61[0:0];
  assign pgassign62[3:3] = BRAM_WEN_A[0:0];
  assign pgassign62[2:2] = BRAM_WEN_A[0:0];
  assign pgassign62[1:1] = BRAM_WEN_A[0:0];
  assign pgassign62[0:0] = BRAM_WEN_A[0:0];
  assign pgassign63[14:14] = 1'b1;
  assign pgassign63[13:0] = BRAM_Addr_B[16:29];
  assign pgassign64[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign64[0:0] = BRAM_Dout_B[7:7];
  assign BRAM_Din_B[7:7] = pgassign65[0:0];
  assign pgassign66[3:3] = BRAM_WEN_B[0:0];
  assign pgassign66[2:2] = BRAM_WEN_B[0:0];
  assign pgassign66[1:1] = BRAM_WEN_B[0:0];
  assign pgassign66[0:0] = BRAM_WEN_B[0:0];
  assign pgassign67[14:14] = 1'b1;
  assign pgassign67[13:0] = BRAM_Addr_A[16:29];
  assign pgassign68[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign68[0:0] = BRAM_Dout_A[8:8];
  assign BRAM_Din_A[8:8] = pgassign69[0:0];
  assign pgassign70[3:3] = BRAM_WEN_A[1:1];
  assign pgassign70[2:2] = BRAM_WEN_A[1:1];
  assign pgassign70[1:1] = BRAM_WEN_A[1:1];
  assign pgassign70[0:0] = BRAM_WEN_A[1:1];
  assign pgassign71[14:14] = 1'b1;
  assign pgassign71[13:0] = BRAM_Addr_B[16:29];
  assign pgassign72[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign72[0:0] = BRAM_Dout_B[8:8];
  assign BRAM_Din_B[8:8] = pgassign73[0:0];
  assign pgassign74[3:3] = BRAM_WEN_B[1:1];
  assign pgassign74[2:2] = BRAM_WEN_B[1:1];
  assign pgassign74[1:1] = BRAM_WEN_B[1:1];
  assign pgassign74[0:0] = BRAM_WEN_B[1:1];
  assign pgassign75[14:14] = 1'b1;
  assign pgassign75[13:0] = BRAM_Addr_A[16:29];
  assign pgassign76[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign76[0:0] = BRAM_Dout_A[9:9];
  assign BRAM_Din_A[9:9] = pgassign77[0:0];
  assign pgassign78[3:3] = BRAM_WEN_A[1:1];
  assign pgassign78[2:2] = BRAM_WEN_A[1:1];
  assign pgassign78[1:1] = BRAM_WEN_A[1:1];
  assign pgassign78[0:0] = BRAM_WEN_A[1:1];
  assign pgassign79[14:14] = 1'b1;
  assign pgassign79[13:0] = BRAM_Addr_B[16:29];
  assign pgassign80[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign80[0:0] = BRAM_Dout_B[9:9];
  assign BRAM_Din_B[9:9] = pgassign81[0:0];
  assign pgassign82[3:3] = BRAM_WEN_B[1:1];
  assign pgassign82[2:2] = BRAM_WEN_B[1:1];
  assign pgassign82[1:1] = BRAM_WEN_B[1:1];
  assign pgassign82[0:0] = BRAM_WEN_B[1:1];
  assign pgassign83[14:14] = 1'b1;
  assign pgassign83[13:0] = BRAM_Addr_A[16:29];
  assign pgassign84[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign84[0:0] = BRAM_Dout_A[10:10];
  assign BRAM_Din_A[10:10] = pgassign85[0:0];
  assign pgassign86[3:3] = BRAM_WEN_A[1:1];
  assign pgassign86[2:2] = BRAM_WEN_A[1:1];
  assign pgassign86[1:1] = BRAM_WEN_A[1:1];
  assign pgassign86[0:0] = BRAM_WEN_A[1:1];
  assign pgassign87[14:14] = 1'b1;
  assign pgassign87[13:0] = BRAM_Addr_B[16:29];
  assign pgassign88[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign88[0:0] = BRAM_Dout_B[10:10];
  assign BRAM_Din_B[10:10] = pgassign89[0:0];
  assign pgassign90[3:3] = BRAM_WEN_B[1:1];
  assign pgassign90[2:2] = BRAM_WEN_B[1:1];
  assign pgassign90[1:1] = BRAM_WEN_B[1:1];
  assign pgassign90[0:0] = BRAM_WEN_B[1:1];
  assign pgassign91[14:14] = 1'b1;
  assign pgassign91[13:0] = BRAM_Addr_A[16:29];
  assign pgassign92[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign92[0:0] = BRAM_Dout_A[11:11];
  assign BRAM_Din_A[11:11] = pgassign93[0:0];
  assign pgassign94[3:3] = BRAM_WEN_A[1:1];
  assign pgassign94[2:2] = BRAM_WEN_A[1:1];
  assign pgassign94[1:1] = BRAM_WEN_A[1:1];
  assign pgassign94[0:0] = BRAM_WEN_A[1:1];
  assign pgassign95[14:14] = 1'b1;
  assign pgassign95[13:0] = BRAM_Addr_B[16:29];
  assign pgassign96[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign96[0:0] = BRAM_Dout_B[11:11];
  assign BRAM_Din_B[11:11] = pgassign97[0:0];
  assign pgassign98[3:3] = BRAM_WEN_B[1:1];
  assign pgassign98[2:2] = BRAM_WEN_B[1:1];
  assign pgassign98[1:1] = BRAM_WEN_B[1:1];
  assign pgassign98[0:0] = BRAM_WEN_B[1:1];
  assign pgassign99[14:14] = 1'b1;
  assign pgassign99[13:0] = BRAM_Addr_A[16:29];
  assign pgassign100[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign100[0:0] = BRAM_Dout_A[12:12];
  assign BRAM_Din_A[12:12] = pgassign101[0:0];
  assign pgassign102[3:3] = BRAM_WEN_A[1:1];
  assign pgassign102[2:2] = BRAM_WEN_A[1:1];
  assign pgassign102[1:1] = BRAM_WEN_A[1:1];
  assign pgassign102[0:0] = BRAM_WEN_A[1:1];
  assign pgassign103[14:14] = 1'b1;
  assign pgassign103[13:0] = BRAM_Addr_B[16:29];
  assign pgassign104[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign104[0:0] = BRAM_Dout_B[12:12];
  assign BRAM_Din_B[12:12] = pgassign105[0:0];
  assign pgassign106[3:3] = BRAM_WEN_B[1:1];
  assign pgassign106[2:2] = BRAM_WEN_B[1:1];
  assign pgassign106[1:1] = BRAM_WEN_B[1:1];
  assign pgassign106[0:0] = BRAM_WEN_B[1:1];
  assign pgassign107[14:14] = 1'b1;
  assign pgassign107[13:0] = BRAM_Addr_A[16:29];
  assign pgassign108[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign108[0:0] = BRAM_Dout_A[13:13];
  assign BRAM_Din_A[13:13] = pgassign109[0:0];
  assign pgassign110[3:3] = BRAM_WEN_A[1:1];
  assign pgassign110[2:2] = BRAM_WEN_A[1:1];
  assign pgassign110[1:1] = BRAM_WEN_A[1:1];
  assign pgassign110[0:0] = BRAM_WEN_A[1:1];
  assign pgassign111[14:14] = 1'b1;
  assign pgassign111[13:0] = BRAM_Addr_B[16:29];
  assign pgassign112[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign112[0:0] = BRAM_Dout_B[13:13];
  assign BRAM_Din_B[13:13] = pgassign113[0:0];
  assign pgassign114[3:3] = BRAM_WEN_B[1:1];
  assign pgassign114[2:2] = BRAM_WEN_B[1:1];
  assign pgassign114[1:1] = BRAM_WEN_B[1:1];
  assign pgassign114[0:0] = BRAM_WEN_B[1:1];
  assign pgassign115[14:14] = 1'b1;
  assign pgassign115[13:0] = BRAM_Addr_A[16:29];
  assign pgassign116[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign116[0:0] = BRAM_Dout_A[14:14];
  assign BRAM_Din_A[14:14] = pgassign117[0:0];
  assign pgassign118[3:3] = BRAM_WEN_A[1:1];
  assign pgassign118[2:2] = BRAM_WEN_A[1:1];
  assign pgassign118[1:1] = BRAM_WEN_A[1:1];
  assign pgassign118[0:0] = BRAM_WEN_A[1:1];
  assign pgassign119[14:14] = 1'b1;
  assign pgassign119[13:0] = BRAM_Addr_B[16:29];
  assign pgassign120[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign120[0:0] = BRAM_Dout_B[14:14];
  assign BRAM_Din_B[14:14] = pgassign121[0:0];
  assign pgassign122[3:3] = BRAM_WEN_B[1:1];
  assign pgassign122[2:2] = BRAM_WEN_B[1:1];
  assign pgassign122[1:1] = BRAM_WEN_B[1:1];
  assign pgassign122[0:0] = BRAM_WEN_B[1:1];
  assign pgassign123[14:14] = 1'b1;
  assign pgassign123[13:0] = BRAM_Addr_A[16:29];
  assign pgassign124[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign124[0:0] = BRAM_Dout_A[15:15];
  assign BRAM_Din_A[15:15] = pgassign125[0:0];
  assign pgassign126[3:3] = BRAM_WEN_A[1:1];
  assign pgassign126[2:2] = BRAM_WEN_A[1:1];
  assign pgassign126[1:1] = BRAM_WEN_A[1:1];
  assign pgassign126[0:0] = BRAM_WEN_A[1:1];
  assign pgassign127[14:14] = 1'b1;
  assign pgassign127[13:0] = BRAM_Addr_B[16:29];
  assign pgassign128[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign128[0:0] = BRAM_Dout_B[15:15];
  assign BRAM_Din_B[15:15] = pgassign129[0:0];
  assign pgassign130[3:3] = BRAM_WEN_B[1:1];
  assign pgassign130[2:2] = BRAM_WEN_B[1:1];
  assign pgassign130[1:1] = BRAM_WEN_B[1:1];
  assign pgassign130[0:0] = BRAM_WEN_B[1:1];
  assign pgassign131[14:14] = 1'b1;
  assign pgassign131[13:0] = BRAM_Addr_A[16:29];
  assign pgassign132[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign132[0:0] = BRAM_Dout_A[16:16];
  assign BRAM_Din_A[16:16] = pgassign133[0:0];
  assign pgassign134[3:3] = BRAM_WEN_A[2:2];
  assign pgassign134[2:2] = BRAM_WEN_A[2:2];
  assign pgassign134[1:1] = BRAM_WEN_A[2:2];
  assign pgassign134[0:0] = BRAM_WEN_A[2:2];
  assign pgassign135[14:14] = 1'b1;
  assign pgassign135[13:0] = BRAM_Addr_B[16:29];
  assign pgassign136[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign136[0:0] = BRAM_Dout_B[16:16];
  assign BRAM_Din_B[16:16] = pgassign137[0:0];
  assign pgassign138[3:3] = BRAM_WEN_B[2:2];
  assign pgassign138[2:2] = BRAM_WEN_B[2:2];
  assign pgassign138[1:1] = BRAM_WEN_B[2:2];
  assign pgassign138[0:0] = BRAM_WEN_B[2:2];
  assign pgassign139[14:14] = 1'b1;
  assign pgassign139[13:0] = BRAM_Addr_A[16:29];
  assign pgassign140[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign140[0:0] = BRAM_Dout_A[17:17];
  assign BRAM_Din_A[17:17] = pgassign141[0:0];
  assign pgassign142[3:3] = BRAM_WEN_A[2:2];
  assign pgassign142[2:2] = BRAM_WEN_A[2:2];
  assign pgassign142[1:1] = BRAM_WEN_A[2:2];
  assign pgassign142[0:0] = BRAM_WEN_A[2:2];
  assign pgassign143[14:14] = 1'b1;
  assign pgassign143[13:0] = BRAM_Addr_B[16:29];
  assign pgassign144[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign144[0:0] = BRAM_Dout_B[17:17];
  assign BRAM_Din_B[17:17] = pgassign145[0:0];
  assign pgassign146[3:3] = BRAM_WEN_B[2:2];
  assign pgassign146[2:2] = BRAM_WEN_B[2:2];
  assign pgassign146[1:1] = BRAM_WEN_B[2:2];
  assign pgassign146[0:0] = BRAM_WEN_B[2:2];
  assign pgassign147[14:14] = 1'b1;
  assign pgassign147[13:0] = BRAM_Addr_A[16:29];
  assign pgassign148[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign148[0:0] = BRAM_Dout_A[18:18];
  assign BRAM_Din_A[18:18] = pgassign149[0:0];
  assign pgassign150[3:3] = BRAM_WEN_A[2:2];
  assign pgassign150[2:2] = BRAM_WEN_A[2:2];
  assign pgassign150[1:1] = BRAM_WEN_A[2:2];
  assign pgassign150[0:0] = BRAM_WEN_A[2:2];
  assign pgassign151[14:14] = 1'b1;
  assign pgassign151[13:0] = BRAM_Addr_B[16:29];
  assign pgassign152[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign152[0:0] = BRAM_Dout_B[18:18];
  assign BRAM_Din_B[18:18] = pgassign153[0:0];
  assign pgassign154[3:3] = BRAM_WEN_B[2:2];
  assign pgassign154[2:2] = BRAM_WEN_B[2:2];
  assign pgassign154[1:1] = BRAM_WEN_B[2:2];
  assign pgassign154[0:0] = BRAM_WEN_B[2:2];
  assign pgassign155[14:14] = 1'b1;
  assign pgassign155[13:0] = BRAM_Addr_A[16:29];
  assign pgassign156[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign156[0:0] = BRAM_Dout_A[19:19];
  assign BRAM_Din_A[19:19] = pgassign157[0:0];
  assign pgassign158[3:3] = BRAM_WEN_A[2:2];
  assign pgassign158[2:2] = BRAM_WEN_A[2:2];
  assign pgassign158[1:1] = BRAM_WEN_A[2:2];
  assign pgassign158[0:0] = BRAM_WEN_A[2:2];
  assign pgassign159[14:14] = 1'b1;
  assign pgassign159[13:0] = BRAM_Addr_B[16:29];
  assign pgassign160[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign160[0:0] = BRAM_Dout_B[19:19];
  assign BRAM_Din_B[19:19] = pgassign161[0:0];
  assign pgassign162[3:3] = BRAM_WEN_B[2:2];
  assign pgassign162[2:2] = BRAM_WEN_B[2:2];
  assign pgassign162[1:1] = BRAM_WEN_B[2:2];
  assign pgassign162[0:0] = BRAM_WEN_B[2:2];
  assign pgassign163[14:14] = 1'b1;
  assign pgassign163[13:0] = BRAM_Addr_A[16:29];
  assign pgassign164[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign164[0:0] = BRAM_Dout_A[20:20];
  assign BRAM_Din_A[20:20] = pgassign165[0:0];
  assign pgassign166[3:3] = BRAM_WEN_A[2:2];
  assign pgassign166[2:2] = BRAM_WEN_A[2:2];
  assign pgassign166[1:1] = BRAM_WEN_A[2:2];
  assign pgassign166[0:0] = BRAM_WEN_A[2:2];
  assign pgassign167[14:14] = 1'b1;
  assign pgassign167[13:0] = BRAM_Addr_B[16:29];
  assign pgassign168[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign168[0:0] = BRAM_Dout_B[20:20];
  assign BRAM_Din_B[20:20] = pgassign169[0:0];
  assign pgassign170[3:3] = BRAM_WEN_B[2:2];
  assign pgassign170[2:2] = BRAM_WEN_B[2:2];
  assign pgassign170[1:1] = BRAM_WEN_B[2:2];
  assign pgassign170[0:0] = BRAM_WEN_B[2:2];
  assign pgassign171[14:14] = 1'b1;
  assign pgassign171[13:0] = BRAM_Addr_A[16:29];
  assign pgassign172[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign172[0:0] = BRAM_Dout_A[21:21];
  assign BRAM_Din_A[21:21] = pgassign173[0:0];
  assign pgassign174[3:3] = BRAM_WEN_A[2:2];
  assign pgassign174[2:2] = BRAM_WEN_A[2:2];
  assign pgassign174[1:1] = BRAM_WEN_A[2:2];
  assign pgassign174[0:0] = BRAM_WEN_A[2:2];
  assign pgassign175[14:14] = 1'b1;
  assign pgassign175[13:0] = BRAM_Addr_B[16:29];
  assign pgassign176[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign176[0:0] = BRAM_Dout_B[21:21];
  assign BRAM_Din_B[21:21] = pgassign177[0:0];
  assign pgassign178[3:3] = BRAM_WEN_B[2:2];
  assign pgassign178[2:2] = BRAM_WEN_B[2:2];
  assign pgassign178[1:1] = BRAM_WEN_B[2:2];
  assign pgassign178[0:0] = BRAM_WEN_B[2:2];
  assign pgassign179[14:14] = 1'b1;
  assign pgassign179[13:0] = BRAM_Addr_A[16:29];
  assign pgassign180[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign180[0:0] = BRAM_Dout_A[22:22];
  assign BRAM_Din_A[22:22] = pgassign181[0:0];
  assign pgassign182[3:3] = BRAM_WEN_A[2:2];
  assign pgassign182[2:2] = BRAM_WEN_A[2:2];
  assign pgassign182[1:1] = BRAM_WEN_A[2:2];
  assign pgassign182[0:0] = BRAM_WEN_A[2:2];
  assign pgassign183[14:14] = 1'b1;
  assign pgassign183[13:0] = BRAM_Addr_B[16:29];
  assign pgassign184[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign184[0:0] = BRAM_Dout_B[22:22];
  assign BRAM_Din_B[22:22] = pgassign185[0:0];
  assign pgassign186[3:3] = BRAM_WEN_B[2:2];
  assign pgassign186[2:2] = BRAM_WEN_B[2:2];
  assign pgassign186[1:1] = BRAM_WEN_B[2:2];
  assign pgassign186[0:0] = BRAM_WEN_B[2:2];
  assign pgassign187[14:14] = 1'b1;
  assign pgassign187[13:0] = BRAM_Addr_A[16:29];
  assign pgassign188[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign188[0:0] = BRAM_Dout_A[23:23];
  assign BRAM_Din_A[23:23] = pgassign189[0:0];
  assign pgassign190[3:3] = BRAM_WEN_A[2:2];
  assign pgassign190[2:2] = BRAM_WEN_A[2:2];
  assign pgassign190[1:1] = BRAM_WEN_A[2:2];
  assign pgassign190[0:0] = BRAM_WEN_A[2:2];
  assign pgassign191[14:14] = 1'b1;
  assign pgassign191[13:0] = BRAM_Addr_B[16:29];
  assign pgassign192[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign192[0:0] = BRAM_Dout_B[23:23];
  assign BRAM_Din_B[23:23] = pgassign193[0:0];
  assign pgassign194[3:3] = BRAM_WEN_B[2:2];
  assign pgassign194[2:2] = BRAM_WEN_B[2:2];
  assign pgassign194[1:1] = BRAM_WEN_B[2:2];
  assign pgassign194[0:0] = BRAM_WEN_B[2:2];
  assign pgassign195[14:14] = 1'b1;
  assign pgassign195[13:0] = BRAM_Addr_A[16:29];
  assign pgassign196[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign196[0:0] = BRAM_Dout_A[24:24];
  assign BRAM_Din_A[24:24] = pgassign197[0:0];
  assign pgassign198[3:3] = BRAM_WEN_A[3:3];
  assign pgassign198[2:2] = BRAM_WEN_A[3:3];
  assign pgassign198[1:1] = BRAM_WEN_A[3:3];
  assign pgassign198[0:0] = BRAM_WEN_A[3:3];
  assign pgassign199[14:14] = 1'b1;
  assign pgassign199[13:0] = BRAM_Addr_B[16:29];
  assign pgassign200[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign200[0:0] = BRAM_Dout_B[24:24];
  assign BRAM_Din_B[24:24] = pgassign201[0:0];
  assign pgassign202[3:3] = BRAM_WEN_B[3:3];
  assign pgassign202[2:2] = BRAM_WEN_B[3:3];
  assign pgassign202[1:1] = BRAM_WEN_B[3:3];
  assign pgassign202[0:0] = BRAM_WEN_B[3:3];
  assign pgassign203[14:14] = 1'b1;
  assign pgassign203[13:0] = BRAM_Addr_A[16:29];
  assign pgassign204[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign204[0:0] = BRAM_Dout_A[25:25];
  assign BRAM_Din_A[25:25] = pgassign205[0:0];
  assign pgassign206[3:3] = BRAM_WEN_A[3:3];
  assign pgassign206[2:2] = BRAM_WEN_A[3:3];
  assign pgassign206[1:1] = BRAM_WEN_A[3:3];
  assign pgassign206[0:0] = BRAM_WEN_A[3:3];
  assign pgassign207[14:14] = 1'b1;
  assign pgassign207[13:0] = BRAM_Addr_B[16:29];
  assign pgassign208[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign208[0:0] = BRAM_Dout_B[25:25];
  assign BRAM_Din_B[25:25] = pgassign209[0:0];
  assign pgassign210[3:3] = BRAM_WEN_B[3:3];
  assign pgassign210[2:2] = BRAM_WEN_B[3:3];
  assign pgassign210[1:1] = BRAM_WEN_B[3:3];
  assign pgassign210[0:0] = BRAM_WEN_B[3:3];
  assign pgassign211[14:14] = 1'b1;
  assign pgassign211[13:0] = BRAM_Addr_A[16:29];
  assign pgassign212[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign212[0:0] = BRAM_Dout_A[26:26];
  assign BRAM_Din_A[26:26] = pgassign213[0:0];
  assign pgassign214[3:3] = BRAM_WEN_A[3:3];
  assign pgassign214[2:2] = BRAM_WEN_A[3:3];
  assign pgassign214[1:1] = BRAM_WEN_A[3:3];
  assign pgassign214[0:0] = BRAM_WEN_A[3:3];
  assign pgassign215[14:14] = 1'b1;
  assign pgassign215[13:0] = BRAM_Addr_B[16:29];
  assign pgassign216[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign216[0:0] = BRAM_Dout_B[26:26];
  assign BRAM_Din_B[26:26] = pgassign217[0:0];
  assign pgassign218[3:3] = BRAM_WEN_B[3:3];
  assign pgassign218[2:2] = BRAM_WEN_B[3:3];
  assign pgassign218[1:1] = BRAM_WEN_B[3:3];
  assign pgassign218[0:0] = BRAM_WEN_B[3:3];
  assign pgassign219[14:14] = 1'b1;
  assign pgassign219[13:0] = BRAM_Addr_A[16:29];
  assign pgassign220[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign220[0:0] = BRAM_Dout_A[27:27];
  assign BRAM_Din_A[27:27] = pgassign221[0:0];
  assign pgassign222[3:3] = BRAM_WEN_A[3:3];
  assign pgassign222[2:2] = BRAM_WEN_A[3:3];
  assign pgassign222[1:1] = BRAM_WEN_A[3:3];
  assign pgassign222[0:0] = BRAM_WEN_A[3:3];
  assign pgassign223[14:14] = 1'b1;
  assign pgassign223[13:0] = BRAM_Addr_B[16:29];
  assign pgassign224[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign224[0:0] = BRAM_Dout_B[27:27];
  assign BRAM_Din_B[27:27] = pgassign225[0:0];
  assign pgassign226[3:3] = BRAM_WEN_B[3:3];
  assign pgassign226[2:2] = BRAM_WEN_B[3:3];
  assign pgassign226[1:1] = BRAM_WEN_B[3:3];
  assign pgassign226[0:0] = BRAM_WEN_B[3:3];
  assign pgassign227[14:14] = 1'b1;
  assign pgassign227[13:0] = BRAM_Addr_A[16:29];
  assign pgassign228[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign228[0:0] = BRAM_Dout_A[28:28];
  assign BRAM_Din_A[28:28] = pgassign229[0:0];
  assign pgassign230[3:3] = BRAM_WEN_A[3:3];
  assign pgassign230[2:2] = BRAM_WEN_A[3:3];
  assign pgassign230[1:1] = BRAM_WEN_A[3:3];
  assign pgassign230[0:0] = BRAM_WEN_A[3:3];
  assign pgassign231[14:14] = 1'b1;
  assign pgassign231[13:0] = BRAM_Addr_B[16:29];
  assign pgassign232[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign232[0:0] = BRAM_Dout_B[28:28];
  assign BRAM_Din_B[28:28] = pgassign233[0:0];
  assign pgassign234[3:3] = BRAM_WEN_B[3:3];
  assign pgassign234[2:2] = BRAM_WEN_B[3:3];
  assign pgassign234[1:1] = BRAM_WEN_B[3:3];
  assign pgassign234[0:0] = BRAM_WEN_B[3:3];
  assign pgassign235[14:14] = 1'b1;
  assign pgassign235[13:0] = BRAM_Addr_A[16:29];
  assign pgassign236[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign236[0:0] = BRAM_Dout_A[29:29];
  assign BRAM_Din_A[29:29] = pgassign237[0:0];
  assign pgassign238[3:3] = BRAM_WEN_A[3:3];
  assign pgassign238[2:2] = BRAM_WEN_A[3:3];
  assign pgassign238[1:1] = BRAM_WEN_A[3:3];
  assign pgassign238[0:0] = BRAM_WEN_A[3:3];
  assign pgassign239[14:14] = 1'b1;
  assign pgassign239[13:0] = BRAM_Addr_B[16:29];
  assign pgassign240[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign240[0:0] = BRAM_Dout_B[29:29];
  assign BRAM_Din_B[29:29] = pgassign241[0:0];
  assign pgassign242[3:3] = BRAM_WEN_B[3:3];
  assign pgassign242[2:2] = BRAM_WEN_B[3:3];
  assign pgassign242[1:1] = BRAM_WEN_B[3:3];
  assign pgassign242[0:0] = BRAM_WEN_B[3:3];
  assign pgassign243[14:14] = 1'b1;
  assign pgassign243[13:0] = BRAM_Addr_A[16:29];
  assign pgassign244[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign244[0:0] = BRAM_Dout_A[30:30];
  assign BRAM_Din_A[30:30] = pgassign245[0:0];
  assign pgassign246[3:3] = BRAM_WEN_A[3:3];
  assign pgassign246[2:2] = BRAM_WEN_A[3:3];
  assign pgassign246[1:1] = BRAM_WEN_A[3:3];
  assign pgassign246[0:0] = BRAM_WEN_A[3:3];
  assign pgassign247[14:14] = 1'b1;
  assign pgassign247[13:0] = BRAM_Addr_B[16:29];
  assign pgassign248[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign248[0:0] = BRAM_Dout_B[30:30];
  assign BRAM_Din_B[30:30] = pgassign249[0:0];
  assign pgassign250[3:3] = BRAM_WEN_B[3:3];
  assign pgassign250[2:2] = BRAM_WEN_B[3:3];
  assign pgassign250[1:1] = BRAM_WEN_B[3:3];
  assign pgassign250[0:0] = BRAM_WEN_B[3:3];
  assign pgassign251[14:14] = 1'b1;
  assign pgassign251[13:0] = BRAM_Addr_A[16:29];
  assign pgassign252[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign252[0:0] = BRAM_Dout_A[31:31];
  assign BRAM_Din_A[31:31] = pgassign253[0:0];
  assign pgassign254[3:3] = BRAM_WEN_A[3:3];
  assign pgassign254[2:2] = BRAM_WEN_A[3:3];
  assign pgassign254[1:1] = BRAM_WEN_A[3:3];
  assign pgassign254[0:0] = BRAM_WEN_A[3:3];
  assign pgassign255[14:14] = 1'b1;
  assign pgassign255[13:0] = BRAM_Addr_B[16:29];
  assign pgassign256[31:1] = 31'b0000000000000000000000000000000;
  assign pgassign256[0:0] = BRAM_Dout_B[31:31];
  assign BRAM_Din_B[31:31] = pgassign257[0:0];
  assign pgassign258[3:3] = BRAM_WEN_B[3:3];
  assign pgassign258[2:2] = BRAM_WEN_B[3:3];
  assign pgassign258[1:1] = BRAM_WEN_B[3:3];
  assign pgassign258[0:0] = BRAM_WEN_B[3:3];
  assign net_gnd0 = 1'b0;
  assign net_gnd4[3:0] = 4'b0000;

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_0.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_0 (
      .ADDRA ( pgassign3 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign4 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign5 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign6 ),
      .ADDRB ( pgassign7 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign8 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign9 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign10 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_1.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_1 (
      .ADDRA ( pgassign11 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign12 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign13 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign14 ),
      .ADDRB ( pgassign15 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign16 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign17 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign18 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_2.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_2 (
      .ADDRA ( pgassign19 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign20 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign21 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign22 ),
      .ADDRB ( pgassign23 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign24 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign25 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign26 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_3.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_3 (
      .ADDRA ( pgassign27 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign28 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign29 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign30 ),
      .ADDRB ( pgassign31 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign32 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign33 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign34 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_4.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_4 (
      .ADDRA ( pgassign35 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign36 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign37 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign38 ),
      .ADDRB ( pgassign39 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign40 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign41 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign42 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_5.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_5 (
      .ADDRA ( pgassign43 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign44 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign45 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign46 ),
      .ADDRB ( pgassign47 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign48 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign49 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign50 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_6.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_6 (
      .ADDRA ( pgassign51 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign52 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign53 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign54 ),
      .ADDRB ( pgassign55 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign56 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign57 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign58 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_7.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_7 (
      .ADDRA ( pgassign59 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign60 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign61 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign62 ),
      .ADDRB ( pgassign63 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign64 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign65 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign66 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_8.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_8 (
      .ADDRA ( pgassign67 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign68 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign69 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign70 ),
      .ADDRB ( pgassign71 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign72 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign73 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign74 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_9.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_9 (
      .ADDRA ( pgassign75 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign76 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign77 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign78 ),
      .ADDRB ( pgassign79 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign80 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign81 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign82 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_10.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_10 (
      .ADDRA ( pgassign83 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign84 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign85 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign86 ),
      .ADDRB ( pgassign87 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign88 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign89 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign90 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_11.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_11 (
      .ADDRA ( pgassign91 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign92 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign93 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign94 ),
      .ADDRB ( pgassign95 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign96 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign97 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign98 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_12.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_12 (
      .ADDRA ( pgassign99 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign100 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign101 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign102 ),
      .ADDRB ( pgassign103 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign104 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign105 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign106 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_13.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_13 (
      .ADDRA ( pgassign107 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign108 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign109 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign110 ),
      .ADDRB ( pgassign111 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign112 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign113 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign114 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_14.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_14 (
      .ADDRA ( pgassign115 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign116 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign117 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign118 ),
      .ADDRB ( pgassign119 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign120 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign121 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign122 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_15.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_15 (
      .ADDRA ( pgassign123 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign124 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign125 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign126 ),
      .ADDRB ( pgassign127 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign128 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign129 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign130 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_16.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_16 (
      .ADDRA ( pgassign131 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign132 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign133 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign134 ),
      .ADDRB ( pgassign135 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign136 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign137 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign138 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_17.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_17 (
      .ADDRA ( pgassign139 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign140 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign141 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign142 ),
      .ADDRB ( pgassign143 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign144 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign145 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign146 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_18.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_18 (
      .ADDRA ( pgassign147 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign148 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign149 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign150 ),
      .ADDRB ( pgassign151 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign152 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign153 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign154 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_19.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_19 (
      .ADDRA ( pgassign155 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign156 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign157 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign158 ),
      .ADDRB ( pgassign159 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign160 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign161 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign162 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_20.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_20 (
      .ADDRA ( pgassign163 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign164 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign165 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign166 ),
      .ADDRB ( pgassign167 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign168 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign169 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign170 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_21.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_21 (
      .ADDRA ( pgassign171 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign172 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign173 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign174 ),
      .ADDRB ( pgassign175 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign176 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign177 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign178 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_22.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_22 (
      .ADDRA ( pgassign179 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign180 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign181 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign182 ),
      .ADDRB ( pgassign183 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign184 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign185 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign186 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_23.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_23 (
      .ADDRA ( pgassign187 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign188 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign189 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign190 ),
      .ADDRB ( pgassign191 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign192 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign193 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign194 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_24.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_24 (
      .ADDRA ( pgassign195 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign196 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign197 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign198 ),
      .ADDRB ( pgassign199 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign200 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign201 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign202 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_25.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_25 (
      .ADDRA ( pgassign203 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign204 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign205 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign206 ),
      .ADDRB ( pgassign207 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign208 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign209 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign210 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_26.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_26 (
      .ADDRA ( pgassign211 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign212 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign213 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign214 ),
      .ADDRB ( pgassign215 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign216 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign217 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign218 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_27.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_27 (
      .ADDRA ( pgassign219 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign220 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign221 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign222 ),
      .ADDRB ( pgassign223 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign224 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign225 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign226 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_28.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_28 (
      .ADDRA ( pgassign227 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign228 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign229 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign230 ),
      .ADDRB ( pgassign231 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign232 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign233 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign234 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_29.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_29 (
      .ADDRA ( pgassign235 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign236 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign237 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign238 ),
      .ADDRB ( pgassign239 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign240 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign241 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign242 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_30.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_30 (
      .ADDRA ( pgassign243 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign244 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign245 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign246 ),
      .ADDRB ( pgassign247 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign248 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign249 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign250 )
    );

  RAMB16
    #(
      .WRITE_MODE_A ( "WRITE_FIRST" ),
      .WRITE_MODE_B ( "WRITE_FIRST" ),
      .INIT_FILE ( "lmb_bram_combined_31.mem" ),
      .READ_WIDTH_A ( 1 ),
      .READ_WIDTH_B ( 1 ),
      .WRITE_WIDTH_A ( 1 ),
      .WRITE_WIDTH_B ( 1 ),
      .RAM_EXTENSION_A ( "NONE" ),
      .RAM_EXTENSION_B ( "NONE" )
    )
    ramb16_31 (
      .ADDRA ( pgassign251 ),
      .CASCADEINA ( net_gnd0 ),
      .CASCADEOUTA (  ),
      .CLKA ( BRAM_Clk_A ),
      .DIA ( pgassign252 ),
      .DIPA ( net_gnd4 ),
      .DOA ( pgassign253 ),
      .DOPA (  ),
      .ENA ( BRAM_EN_A ),
      .REGCEA ( net_gnd0 ),
      .SSRA ( BRAM_Rst_A ),
      .WEA ( pgassign254 ),
      .ADDRB ( pgassign255 ),
      .CASCADEINB ( net_gnd0 ),
      .CASCADEOUTB (  ),
      .CLKB ( BRAM_Clk_B ),
      .DIB ( pgassign256 ),
      .DIPB ( net_gnd4 ),
      .DOB ( pgassign257 ),
      .DOPB (  ),
      .ENB ( BRAM_EN_B ),
      .REGCEB ( net_gnd0 ),
      .SSRB ( BRAM_Rst_B ),
      .WEB ( pgassign258 )
    );

endmodule

