//-----------------------------------------------------------------------------
// microblaze.v
//-----------------------------------------------------------------------------

`timescale 1 ps / 100 fs

`uselib lib=unisims_ver

module microblaze
  (
    fpga_0_RS232_RX_pin,
    fpga_0_RS232_TX_pin,
    fpga_0_clk_1_sys_clk_pin,
    fpga_0_rst_1_sys_rst_pin,
    plb_dac_0_S_Data_pin,
    plb_dac_0_S_DCLKIO_pin,
    plb_dac_0_S_Clkout_pin,
    plb_dac_0_S_PinMD_pin,
    plb_dac_0_S_ClkMD_pin,
    plb_dac_0_S_Format_pin,
    plb_dac_0_S_PWRDN_pin
  );
  input fpga_0_RS232_RX_pin;
  output fpga_0_RS232_TX_pin;
  input fpga_0_clk_1_sys_clk_pin;
  input fpga_0_rst_1_sys_rst_pin;
  output [0:9] plb_dac_0_S_Data_pin;
  output plb_dac_0_S_DCLKIO_pin;
  output plb_dac_0_S_Clkout_pin;
  output plb_dac_0_S_PinMD_pin;
  output plb_dac_0_S_ClkMD_pin;
  output plb_dac_0_S_Format_pin;
  output plb_dac_0_S_PWRDN_pin;

  // Internal signals

  wire CLK_S;
  wire Dcm_all_locked;
  wire Debug_SYS_Rst;
  wire Ext_BRK;
  wire Ext_NM_BRK;
  wire [0:0] RS232_Interrupt;
  wire clk_50_0000MHz;
  wire [0:31] dlmb_LMB_ABus;
  wire dlmb_LMB_AddrStrobe;
  wire [0:3] dlmb_LMB_BE;
  wire dlmb_LMB_CE;
  wire [0:31] dlmb_LMB_ReadDBus;
  wire dlmb_LMB_ReadStrobe;
  wire dlmb_LMB_Ready;
  wire dlmb_LMB_Rst;
  wire dlmb_LMB_UE;
  wire dlmb_LMB_Wait;
  wire [0:31] dlmb_LMB_WriteDBus;
  wire dlmb_LMB_WriteStrobe;
  wire [0:31] dlmb_M_ABus;
  wire dlmb_M_AddrStrobe;
  wire [0:3] dlmb_M_BE;
  wire [0:31] dlmb_M_DBus;
  wire dlmb_M_ReadStrobe;
  wire dlmb_M_WriteStrobe;
  wire [0:0] dlmb_Sl_CE;
  wire [0:31] dlmb_Sl_DBus;
  wire [0:0] dlmb_Sl_Ready;
  wire [0:0] dlmb_Sl_UE;
  wire [0:0] dlmb_Sl_Wait;
  wire [0:31] dlmb_port_BRAM_Addr;
  wire dlmb_port_BRAM_Clk;
  wire [0:31] dlmb_port_BRAM_Din;
  wire [0:31] dlmb_port_BRAM_Dout;
  wire dlmb_port_BRAM_EN;
  wire dlmb_port_BRAM_Rst;
  wire [0:3] dlmb_port_BRAM_WEN;
  wire [0:31] ilmb_LMB_ABus;
  wire ilmb_LMB_AddrStrobe;
  wire [0:3] ilmb_LMB_BE;
  wire ilmb_LMB_CE;
  wire [0:31] ilmb_LMB_ReadDBus;
  wire ilmb_LMB_ReadStrobe;
  wire ilmb_LMB_Ready;
  wire ilmb_LMB_Rst;
  wire ilmb_LMB_UE;
  wire ilmb_LMB_Wait;
  wire [0:31] ilmb_LMB_WriteDBus;
  wire ilmb_LMB_WriteStrobe;
  wire [0:31] ilmb_M_ABus;
  wire ilmb_M_AddrStrobe;
  wire ilmb_M_ReadStrobe;
  wire [0:0] ilmb_Sl_CE;
  wire [0:31] ilmb_Sl_DBus;
  wire [0:0] ilmb_Sl_Ready;
  wire [0:0] ilmb_Sl_UE;
  wire [0:0] ilmb_Sl_Wait;
  wire [0:31] ilmb_cntlr_BRAM_PORT_BRAM_Addr;
  wire ilmb_cntlr_BRAM_PORT_BRAM_Clk;
  wire [0:31] ilmb_cntlr_BRAM_PORT_BRAM_Din;
  wire [0:31] ilmb_cntlr_BRAM_PORT_BRAM_Dout;
  wire ilmb_cntlr_BRAM_PORT_BRAM_EN;
  wire ilmb_cntlr_BRAM_PORT_BRAM_Rst;
  wire [0:3] ilmb_cntlr_BRAM_PORT_BRAM_WEN;
  wire [0:1] mb_plb_M_ABort;
  wire [0:63] mb_plb_M_ABus;
  wire [0:7] mb_plb_M_BE;
  wire [0:3] mb_plb_M_MSize;
  wire [0:1] mb_plb_M_RNW;
  wire [0:31] mb_plb_M_TAttribute;
  wire [0:63] mb_plb_M_UABus;
  wire [0:1] mb_plb_M_busLock;
  wire [0:1] mb_plb_M_lockErr;
  wire [0:3] mb_plb_M_priority;
  wire [0:1] mb_plb_M_rdBurst;
  wire [0:1] mb_plb_M_request;
  wire [0:7] mb_plb_M_size;
  wire [0:5] mb_plb_M_type;
  wire [0:1] mb_plb_M_wrBurst;
  wire [0:63] mb_plb_M_wrDBus;
  wire [0:31] mb_plb_PLB_ABus;
  wire [0:3] mb_plb_PLB_BE;
  wire [0:1] mb_plb_PLB_MAddrAck;
  wire [0:1] mb_plb_PLB_MBusy;
  wire [0:1] mb_plb_PLB_MIRQ;
  wire [0:1] mb_plb_PLB_MRdBTerm;
  wire [0:1] mb_plb_PLB_MRdDAck;
  wire [0:63] mb_plb_PLB_MRdDBus;
  wire [0:1] mb_plb_PLB_MRdErr;
  wire [0:7] mb_plb_PLB_MRdWdAddr;
  wire [0:1] mb_plb_PLB_MRearbitrate;
  wire [0:3] mb_plb_PLB_MSSize;
  wire [0:1] mb_plb_PLB_MSize;
  wire [0:1] mb_plb_PLB_MTimeout;
  wire [0:1] mb_plb_PLB_MWrBTerm;
  wire [0:1] mb_plb_PLB_MWrDAck;
  wire [0:1] mb_plb_PLB_MWrErr;
  wire mb_plb_PLB_PAValid;
  wire mb_plb_PLB_RNW;
  wire mb_plb_PLB_SAValid;
  wire [0:15] mb_plb_PLB_TAttribute;
  wire [0:31] mb_plb_PLB_UABus;
  wire mb_plb_PLB_abort;
  wire mb_plb_PLB_busLock;
  wire mb_plb_PLB_lockErr;
  wire [0:0] mb_plb_PLB_masterID;
  wire mb_plb_PLB_rdBurst;
  wire [0:1] mb_plb_PLB_rdPendPri;
  wire mb_plb_PLB_rdPendReq;
  wire [0:3] mb_plb_PLB_rdPrim;
  wire [0:1] mb_plb_PLB_reqPri;
  wire [0:3] mb_plb_PLB_size;
  wire [0:2] mb_plb_PLB_type;
  wire mb_plb_PLB_wrBurst;
  wire [0:31] mb_plb_PLB_wrDBus;
  wire [0:1] mb_plb_PLB_wrPendPri;
  wire mb_plb_PLB_wrPendReq;
  wire [0:3] mb_plb_PLB_wrPrim;
  wire [0:3] mb_plb_SPLB_Rst;
  wire [0:7] mb_plb_Sl_MBusy;
  wire [0:7] mb_plb_Sl_MIRQ;
  wire [0:7] mb_plb_Sl_MRdErr;
  wire [0:7] mb_plb_Sl_MWrErr;
  wire [0:7] mb_plb_Sl_SSize;
  wire [0:3] mb_plb_Sl_addrAck;
  wire [0:3] mb_plb_Sl_rdBTerm;
  wire [0:3] mb_plb_Sl_rdComp;
  wire [0:3] mb_plb_Sl_rdDAck;
  wire [0:127] mb_plb_Sl_rdDBus;
  wire [0:15] mb_plb_Sl_rdWdAddr;
  wire [0:3] mb_plb_Sl_rearbitrate;
  wire [0:3] mb_plb_Sl_wait;
  wire [0:3] mb_plb_Sl_wrBTerm;
  wire [0:3] mb_plb_Sl_wrComp;
  wire [0:3] mb_plb_Sl_wrDAck;
  wire mb_reset;
  wire microblaze_0_Interrupt;
  wire microblaze_0_mdm_bus_Dbg_Capture;
  wire microblaze_0_mdm_bus_Dbg_Clk;
  wire [0:7] microblaze_0_mdm_bus_Dbg_Reg_En;
  wire microblaze_0_mdm_bus_Dbg_Shift;
  wire microblaze_0_mdm_bus_Dbg_TDI;
  wire microblaze_0_mdm_bus_Dbg_TDO;
  wire microblaze_0_mdm_bus_Dbg_Update;
  wire microblaze_0_mdm_bus_Debug_Rst;
  wire net_gnd0;
  wire [0:0] net_gnd1;
  wire [0:1] net_gnd2;
  wire [2:0] net_gnd3;
  wire [0:3] net_gnd4;
  wire [0:9] net_gnd10;
  wire [0:15] net_gnd16;
  wire [0:31] net_gnd32;
  wire [0:4095] net_gnd4096;
  wire net_vcc0;
  wire plb_dac_0_S_ClkMD;
  wire plb_dac_0_S_Clkout;
  wire plb_dac_0_S_DCLKIO;
  wire [0:9] plb_dac_0_S_Data;
  wire plb_dac_0_S_Format;
  wire plb_dac_0_S_PWRDN;
  wire plb_dac_0_S_PinMD;
  wire [0:0] sys_bus_reset;
  wire sys_rst_s;

  // Internal assignments

  assign CLK_S = fpga_0_clk_1_sys_clk_pin;
  assign sys_rst_s = fpga_0_rst_1_sys_rst_pin;
  assign plb_dac_0_S_Data_pin = plb_dac_0_S_Data;
  assign plb_dac_0_S_DCLKIO_pin = plb_dac_0_S_DCLKIO;
  assign plb_dac_0_S_Clkout_pin = plb_dac_0_S_Clkout;
  assign plb_dac_0_S_PinMD_pin = plb_dac_0_S_PinMD;
  assign plb_dac_0_S_ClkMD_pin = plb_dac_0_S_ClkMD;
  assign plb_dac_0_S_Format_pin = plb_dac_0_S_Format;
  assign plb_dac_0_S_PWRDN_pin = plb_dac_0_S_PWRDN;
  assign net_gnd0 = 1'b0;
  assign net_gnd1[0:0] = 1'b0;
  assign net_gnd10[0:9] = 10'b0000000000;
  assign net_gnd16[0:15] = 16'b0000000000000000;
  assign net_gnd2[0:1] = 2'b00;
  assign net_gnd3[2:0] = 3'b000;
  assign net_gnd32[0:31] = 32'b00000000000000000000000000000000;
  assign net_gnd4[0:3] = 4'b0000;
  assign net_gnd4096[0:4095] = 4096'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign net_vcc0 = 1'b1;

  microblaze_microblaze_0_wrapper
    microblaze_0 (
      .CLK ( clk_50_0000MHz ),
      .RESET ( dlmb_LMB_Rst ),
      .MB_RESET ( mb_reset ),
      .INTERRUPT ( microblaze_0_Interrupt ),
      .INTERRUPT_ADDRESS ( net_gnd32 ),
      .INTERRUPT_ACK (  ),
      .EXT_BRK ( Ext_BRK ),
      .EXT_NM_BRK ( Ext_NM_BRK ),
      .DBG_STOP ( net_gnd0 ),
      .MB_Halted (  ),
      .MB_Error (  ),
      .WAKEUP ( net_gnd2 ),
      .SLEEP (  ),
      .DBG_WAKEUP (  ),
      .LOCKSTEP_MASTER_OUT (  ),
      .LOCKSTEP_SLAVE_IN ( net_gnd4096 ),
      .LOCKSTEP_OUT (  ),
      .INSTR ( ilmb_LMB_ReadDBus ),
      .IREADY ( ilmb_LMB_Ready ),
      .IWAIT ( ilmb_LMB_Wait ),
      .ICE ( ilmb_LMB_CE ),
      .IUE ( ilmb_LMB_UE ),
      .INSTR_ADDR ( ilmb_M_ABus ),
      .IFETCH ( ilmb_M_ReadStrobe ),
      .I_AS ( ilmb_M_AddrStrobe ),
      .IPLB_M_ABort ( mb_plb_M_ABort[1] ),
      .IPLB_M_ABus ( mb_plb_M_ABus[32:63] ),
      .IPLB_M_UABus ( mb_plb_M_UABus[32:63] ),
      .IPLB_M_BE ( mb_plb_M_BE[4:7] ),
      .IPLB_M_busLock ( mb_plb_M_busLock[1] ),
      .IPLB_M_lockErr ( mb_plb_M_lockErr[1] ),
      .IPLB_M_MSize ( mb_plb_M_MSize[2:3] ),
      .IPLB_M_priority ( mb_plb_M_priority[2:3] ),
      .IPLB_M_rdBurst ( mb_plb_M_rdBurst[1] ),
      .IPLB_M_request ( mb_plb_M_request[1] ),
      .IPLB_M_RNW ( mb_plb_M_RNW[1] ),
      .IPLB_M_size ( mb_plb_M_size[4:7] ),
      .IPLB_M_TAttribute ( mb_plb_M_TAttribute[16:31] ),
      .IPLB_M_type ( mb_plb_M_type[3:5] ),
      .IPLB_M_wrBurst ( mb_plb_M_wrBurst[1] ),
      .IPLB_M_wrDBus ( mb_plb_M_wrDBus[32:63] ),
      .IPLB_MBusy ( mb_plb_PLB_MBusy[1] ),
      .IPLB_MRdErr ( mb_plb_PLB_MRdErr[1] ),
      .IPLB_MWrErr ( mb_plb_PLB_MWrErr[1] ),
      .IPLB_MIRQ ( mb_plb_PLB_MIRQ[1] ),
      .IPLB_MWrBTerm ( mb_plb_PLB_MWrBTerm[1] ),
      .IPLB_MWrDAck ( mb_plb_PLB_MWrDAck[1] ),
      .IPLB_MAddrAck ( mb_plb_PLB_MAddrAck[1] ),
      .IPLB_MRdBTerm ( mb_plb_PLB_MRdBTerm[1] ),
      .IPLB_MRdDAck ( mb_plb_PLB_MRdDAck[1] ),
      .IPLB_MRdDBus ( mb_plb_PLB_MRdDBus[32:63] ),
      .IPLB_MRdWdAddr ( mb_plb_PLB_MRdWdAddr[4:7] ),
      .IPLB_MRearbitrate ( mb_plb_PLB_MRearbitrate[1] ),
      .IPLB_MSSize ( mb_plb_PLB_MSSize[2:3] ),
      .IPLB_MTimeout ( mb_plb_PLB_MTimeout[1] ),
      .DATA_READ ( dlmb_LMB_ReadDBus ),
      .DREADY ( dlmb_LMB_Ready ),
      .DWAIT ( dlmb_LMB_Wait ),
      .DCE ( dlmb_LMB_CE ),
      .DUE ( dlmb_LMB_UE ),
      .DATA_WRITE ( dlmb_M_DBus ),
      .DATA_ADDR ( dlmb_M_ABus ),
      .D_AS ( dlmb_M_AddrStrobe ),
      .READ_STROBE ( dlmb_M_ReadStrobe ),
      .WRITE_STROBE ( dlmb_M_WriteStrobe ),
      .BYTE_ENABLE ( dlmb_M_BE ),
      .DPLB_M_ABort ( mb_plb_M_ABort[0] ),
      .DPLB_M_ABus ( mb_plb_M_ABus[0:31] ),
      .DPLB_M_UABus ( mb_plb_M_UABus[0:31] ),
      .DPLB_M_BE ( mb_plb_M_BE[0:3] ),
      .DPLB_M_busLock ( mb_plb_M_busLock[0] ),
      .DPLB_M_lockErr ( mb_plb_M_lockErr[0] ),
      .DPLB_M_MSize ( mb_plb_M_MSize[0:1] ),
      .DPLB_M_priority ( mb_plb_M_priority[0:1] ),
      .DPLB_M_rdBurst ( mb_plb_M_rdBurst[0] ),
      .DPLB_M_request ( mb_plb_M_request[0] ),
      .DPLB_M_RNW ( mb_plb_M_RNW[0] ),
      .DPLB_M_size ( mb_plb_M_size[0:3] ),
      .DPLB_M_TAttribute ( mb_plb_M_TAttribute[0:15] ),
      .DPLB_M_type ( mb_plb_M_type[0:2] ),
      .DPLB_M_wrBurst ( mb_plb_M_wrBurst[0] ),
      .DPLB_M_wrDBus ( mb_plb_M_wrDBus[0:31] ),
      .DPLB_MBusy ( mb_plb_PLB_MBusy[0] ),
      .DPLB_MRdErr ( mb_plb_PLB_MRdErr[0] ),
      .DPLB_MWrErr ( mb_plb_PLB_MWrErr[0] ),
      .DPLB_MIRQ ( mb_plb_PLB_MIRQ[0] ),
      .DPLB_MWrBTerm ( mb_plb_PLB_MWrBTerm[0] ),
      .DPLB_MWrDAck ( mb_plb_PLB_MWrDAck[0] ),
      .DPLB_MAddrAck ( mb_plb_PLB_MAddrAck[0] ),
      .DPLB_MRdBTerm ( mb_plb_PLB_MRdBTerm[0] ),
      .DPLB_MRdDAck ( mb_plb_PLB_MRdDAck[0] ),
      .DPLB_MRdDBus ( mb_plb_PLB_MRdDBus[0:31] ),
      .DPLB_MRdWdAddr ( mb_plb_PLB_MRdWdAddr[0:3] ),
      .DPLB_MRearbitrate ( mb_plb_PLB_MRearbitrate[0] ),
      .DPLB_MSSize ( mb_plb_PLB_MSSize[0:1] ),
      .DPLB_MTimeout ( mb_plb_PLB_MTimeout[0] ),
      .M_AXI_IP_AWID (  ),
      .M_AXI_IP_AWADDR (  ),
      .M_AXI_IP_AWLEN (  ),
      .M_AXI_IP_AWSIZE (  ),
      .M_AXI_IP_AWBURST (  ),
      .M_AXI_IP_AWLOCK (  ),
      .M_AXI_IP_AWCACHE (  ),
      .M_AXI_IP_AWPROT (  ),
      .M_AXI_IP_AWQOS (  ),
      .M_AXI_IP_AWVALID (  ),
      .M_AXI_IP_AWREADY ( net_gnd0 ),
      .M_AXI_IP_WDATA (  ),
      .M_AXI_IP_WSTRB (  ),
      .M_AXI_IP_WLAST (  ),
      .M_AXI_IP_WVALID (  ),
      .M_AXI_IP_WREADY ( net_gnd0 ),
      .M_AXI_IP_BID ( net_gnd1[0:0] ),
      .M_AXI_IP_BRESP ( net_gnd2[0:1] ),
      .M_AXI_IP_BVALID ( net_gnd0 ),
      .M_AXI_IP_BREADY (  ),
      .M_AXI_IP_ARID (  ),
      .M_AXI_IP_ARADDR (  ),
      .M_AXI_IP_ARLEN (  ),
      .M_AXI_IP_ARSIZE (  ),
      .M_AXI_IP_ARBURST (  ),
      .M_AXI_IP_ARLOCK (  ),
      .M_AXI_IP_ARCACHE (  ),
      .M_AXI_IP_ARPROT (  ),
      .M_AXI_IP_ARQOS (  ),
      .M_AXI_IP_ARVALID (  ),
      .M_AXI_IP_ARREADY ( net_gnd0 ),
      .M_AXI_IP_RID ( net_gnd1[0:0] ),
      .M_AXI_IP_RDATA ( net_gnd32[0:31] ),
      .M_AXI_IP_RRESP ( net_gnd2[0:1] ),
      .M_AXI_IP_RLAST ( net_gnd0 ),
      .M_AXI_IP_RVALID ( net_gnd0 ),
      .M_AXI_IP_RREADY (  ),
      .M_AXI_DP_AWID (  ),
      .M_AXI_DP_AWADDR (  ),
      .M_AXI_DP_AWLEN (  ),
      .M_AXI_DP_AWSIZE (  ),
      .M_AXI_DP_AWBURST (  ),
      .M_AXI_DP_AWLOCK (  ),
      .M_AXI_DP_AWCACHE (  ),
      .M_AXI_DP_AWPROT (  ),
      .M_AXI_DP_AWQOS (  ),
      .M_AXI_DP_AWVALID (  ),
      .M_AXI_DP_AWREADY ( net_gnd0 ),
      .M_AXI_DP_WDATA (  ),
      .M_AXI_DP_WSTRB (  ),
      .M_AXI_DP_WLAST (  ),
      .M_AXI_DP_WVALID (  ),
      .M_AXI_DP_WREADY ( net_gnd0 ),
      .M_AXI_DP_BID ( net_gnd1[0:0] ),
      .M_AXI_DP_BRESP ( net_gnd2[0:1] ),
      .M_AXI_DP_BVALID ( net_gnd0 ),
      .M_AXI_DP_BREADY (  ),
      .M_AXI_DP_ARID (  ),
      .M_AXI_DP_ARADDR (  ),
      .M_AXI_DP_ARLEN (  ),
      .M_AXI_DP_ARSIZE (  ),
      .M_AXI_DP_ARBURST (  ),
      .M_AXI_DP_ARLOCK (  ),
      .M_AXI_DP_ARCACHE (  ),
      .M_AXI_DP_ARPROT (  ),
      .M_AXI_DP_ARQOS (  ),
      .M_AXI_DP_ARVALID (  ),
      .M_AXI_DP_ARREADY ( net_gnd0 ),
      .M_AXI_DP_RID ( net_gnd1[0:0] ),
      .M_AXI_DP_RDATA ( net_gnd32[0:31] ),
      .M_AXI_DP_RRESP ( net_gnd2[0:1] ),
      .M_AXI_DP_RLAST ( net_gnd0 ),
      .M_AXI_DP_RVALID ( net_gnd0 ),
      .M_AXI_DP_RREADY (  ),
      .M_AXI_IC_AWID (  ),
      .M_AXI_IC_AWADDR (  ),
      .M_AXI_IC_AWLEN (  ),
      .M_AXI_IC_AWSIZE (  ),
      .M_AXI_IC_AWBURST (  ),
      .M_AXI_IC_AWLOCK (  ),
      .M_AXI_IC_AWCACHE (  ),
      .M_AXI_IC_AWPROT (  ),
      .M_AXI_IC_AWQOS (  ),
      .M_AXI_IC_AWVALID (  ),
      .M_AXI_IC_AWREADY ( net_gnd0 ),
      .M_AXI_IC_AWUSER (  ),
      .M_AXI_IC_AWDOMAIN (  ),
      .M_AXI_IC_AWSNOOP (  ),
      .M_AXI_IC_AWBAR (  ),
      .M_AXI_IC_WDATA (  ),
      .M_AXI_IC_WSTRB (  ),
      .M_AXI_IC_WLAST (  ),
      .M_AXI_IC_WVALID (  ),
      .M_AXI_IC_WREADY ( net_gnd0 ),
      .M_AXI_IC_WUSER (  ),
      .M_AXI_IC_BID ( net_gnd1[0:0] ),
      .M_AXI_IC_BRESP ( net_gnd2[0:1] ),
      .M_AXI_IC_BVALID ( net_gnd0 ),
      .M_AXI_IC_BREADY (  ),
      .M_AXI_IC_BUSER ( net_gnd1[0:0] ),
      .M_AXI_IC_WACK (  ),
      .M_AXI_IC_ARID (  ),
      .M_AXI_IC_ARADDR (  ),
      .M_AXI_IC_ARLEN (  ),
      .M_AXI_IC_ARSIZE (  ),
      .M_AXI_IC_ARBURST (  ),
      .M_AXI_IC_ARLOCK (  ),
      .M_AXI_IC_ARCACHE (  ),
      .M_AXI_IC_ARPROT (  ),
      .M_AXI_IC_ARQOS (  ),
      .M_AXI_IC_ARVALID (  ),
      .M_AXI_IC_ARREADY ( net_gnd0 ),
      .M_AXI_IC_ARUSER (  ),
      .M_AXI_IC_ARDOMAIN (  ),
      .M_AXI_IC_ARSNOOP (  ),
      .M_AXI_IC_ARBAR (  ),
      .M_AXI_IC_RID ( net_gnd1[0:0] ),
      .M_AXI_IC_RDATA ( net_gnd32[0:31] ),
      .M_AXI_IC_RRESP ( net_gnd2[0:1] ),
      .M_AXI_IC_RLAST ( net_gnd0 ),
      .M_AXI_IC_RVALID ( net_gnd0 ),
      .M_AXI_IC_RREADY (  ),
      .M_AXI_IC_RUSER ( net_gnd1[0:0] ),
      .M_AXI_IC_RACK (  ),
      .M_AXI_IC_ACVALID ( net_gnd0 ),
      .M_AXI_IC_ACADDR ( net_gnd32[0:31] ),
      .M_AXI_IC_ACSNOOP ( net_gnd4[0:3] ),
      .M_AXI_IC_ACPROT ( net_gnd3 ),
      .M_AXI_IC_ACREADY (  ),
      .M_AXI_IC_CRREADY ( net_gnd0 ),
      .M_AXI_IC_CRVALID (  ),
      .M_AXI_IC_CRRESP (  ),
      .M_AXI_IC_CDVALID (  ),
      .M_AXI_IC_CDREADY ( net_gnd0 ),
      .M_AXI_IC_CDDATA (  ),
      .M_AXI_IC_CDLAST (  ),
      .M_AXI_DC_AWID (  ),
      .M_AXI_DC_AWADDR (  ),
      .M_AXI_DC_AWLEN (  ),
      .M_AXI_DC_AWSIZE (  ),
      .M_AXI_DC_AWBURST (  ),
      .M_AXI_DC_AWLOCK (  ),
      .M_AXI_DC_AWCACHE (  ),
      .M_AXI_DC_AWPROT (  ),
      .M_AXI_DC_AWQOS (  ),
      .M_AXI_DC_AWVALID (  ),
      .M_AXI_DC_AWREADY ( net_gnd0 ),
      .M_AXI_DC_AWUSER (  ),
      .M_AXI_DC_AWDOMAIN (  ),
      .M_AXI_DC_AWSNOOP (  ),
      .M_AXI_DC_AWBAR (  ),
      .M_AXI_DC_WDATA (  ),
      .M_AXI_DC_WSTRB (  ),
      .M_AXI_DC_WLAST (  ),
      .M_AXI_DC_WVALID (  ),
      .M_AXI_DC_WREADY ( net_gnd0 ),
      .M_AXI_DC_WUSER (  ),
      .M_AXI_DC_BID ( net_gnd1[0:0] ),
      .M_AXI_DC_BRESP ( net_gnd2[0:1] ),
      .M_AXI_DC_BVALID ( net_gnd0 ),
      .M_AXI_DC_BREADY (  ),
      .M_AXI_DC_BUSER ( net_gnd1[0:0] ),
      .M_AXI_DC_WACK (  ),
      .M_AXI_DC_ARID (  ),
      .M_AXI_DC_ARADDR (  ),
      .M_AXI_DC_ARLEN (  ),
      .M_AXI_DC_ARSIZE (  ),
      .M_AXI_DC_ARBURST (  ),
      .M_AXI_DC_ARLOCK (  ),
      .M_AXI_DC_ARCACHE (  ),
      .M_AXI_DC_ARPROT (  ),
      .M_AXI_DC_ARQOS (  ),
      .M_AXI_DC_ARVALID (  ),
      .M_AXI_DC_ARREADY ( net_gnd0 ),
      .M_AXI_DC_ARUSER (  ),
      .M_AXI_DC_ARDOMAIN (  ),
      .M_AXI_DC_ARSNOOP (  ),
      .M_AXI_DC_ARBAR (  ),
      .M_AXI_DC_RID ( net_gnd1[0:0] ),
      .M_AXI_DC_RDATA ( net_gnd32[0:31] ),
      .M_AXI_DC_RRESP ( net_gnd2[0:1] ),
      .M_AXI_DC_RLAST ( net_gnd0 ),
      .M_AXI_DC_RVALID ( net_gnd0 ),
      .M_AXI_DC_RREADY (  ),
      .M_AXI_DC_RUSER ( net_gnd1[0:0] ),
      .M_AXI_DC_RACK (  ),
      .M_AXI_DC_ACVALID ( net_gnd0 ),
      .M_AXI_DC_ACADDR ( net_gnd32[0:31] ),
      .M_AXI_DC_ACSNOOP ( net_gnd4[0:3] ),
      .M_AXI_DC_ACPROT ( net_gnd3 ),
      .M_AXI_DC_ACREADY (  ),
      .M_AXI_DC_CRREADY ( net_gnd0 ),
      .M_AXI_DC_CRVALID (  ),
      .M_AXI_DC_CRRESP (  ),
      .M_AXI_DC_CDVALID (  ),
      .M_AXI_DC_CDREADY ( net_gnd0 ),
      .M_AXI_DC_CDDATA (  ),
      .M_AXI_DC_CDLAST (  ),
      .DBG_CLK ( microblaze_0_mdm_bus_Dbg_Clk ),
      .DBG_TDI ( microblaze_0_mdm_bus_Dbg_TDI ),
      .DBG_TDO ( microblaze_0_mdm_bus_Dbg_TDO ),
      .DBG_REG_EN ( microblaze_0_mdm_bus_Dbg_Reg_En ),
      .DBG_SHIFT ( microblaze_0_mdm_bus_Dbg_Shift ),
      .DBG_CAPTURE ( microblaze_0_mdm_bus_Dbg_Capture ),
      .DBG_UPDATE ( microblaze_0_mdm_bus_Dbg_Update ),
      .DEBUG_RST ( microblaze_0_mdm_bus_Debug_Rst ),
      .Trace_Instruction (  ),
      .Trace_Valid_Instr (  ),
      .Trace_PC (  ),
      .Trace_Reg_Write (  ),
      .Trace_Reg_Addr (  ),
      .Trace_MSR_Reg (  ),
      .Trace_PID_Reg (  ),
      .Trace_New_Reg_Value (  ),
      .Trace_Exception_Taken (  ),
      .Trace_Exception_Kind (  ),
      .Trace_Jump_Taken (  ),
      .Trace_Delay_Slot (  ),
      .Trace_Data_Address (  ),
      .Trace_Data_Access (  ),
      .Trace_Data_Read (  ),
      .Trace_Data_Write (  ),
      .Trace_Data_Write_Value (  ),
      .Trace_Data_Byte_Enable (  ),
      .Trace_DCache_Req (  ),
      .Trace_DCache_Hit (  ),
      .Trace_DCache_Rdy (  ),
      .Trace_DCache_Read (  ),
      .Trace_ICache_Req (  ),
      .Trace_ICache_Hit (  ),
      .Trace_ICache_Rdy (  ),
      .Trace_OF_PipeRun (  ),
      .Trace_EX_PipeRun (  ),
      .Trace_MEM_PipeRun (  ),
      .Trace_MB_Halted (  ),
      .Trace_Jump_Hit (  ),
      .FSL0_S_CLK (  ),
      .FSL0_S_READ (  ),
      .FSL0_S_DATA ( net_gnd32 ),
      .FSL0_S_CONTROL ( net_gnd0 ),
      .FSL0_S_EXISTS ( net_gnd0 ),
      .FSL0_M_CLK (  ),
      .FSL0_M_WRITE (  ),
      .FSL0_M_DATA (  ),
      .FSL0_M_CONTROL (  ),
      .FSL0_M_FULL ( net_gnd0 ),
      .FSL1_S_CLK (  ),
      .FSL1_S_READ (  ),
      .FSL1_S_DATA ( net_gnd32 ),
      .FSL1_S_CONTROL ( net_gnd0 ),
      .FSL1_S_EXISTS ( net_gnd0 ),
      .FSL1_M_CLK (  ),
      .FSL1_M_WRITE (  ),
      .FSL1_M_DATA (  ),
      .FSL1_M_CONTROL (  ),
      .FSL1_M_FULL ( net_gnd0 ),
      .FSL2_S_CLK (  ),
      .FSL2_S_READ (  ),
      .FSL2_S_DATA ( net_gnd32 ),
      .FSL2_S_CONTROL ( net_gnd0 ),
      .FSL2_S_EXISTS ( net_gnd0 ),
      .FSL2_M_CLK (  ),
      .FSL2_M_WRITE (  ),
      .FSL2_M_DATA (  ),
      .FSL2_M_CONTROL (  ),
      .FSL2_M_FULL ( net_gnd0 ),
      .FSL3_S_CLK (  ),
      .FSL3_S_READ (  ),
      .FSL3_S_DATA ( net_gnd32 ),
      .FSL3_S_CONTROL ( net_gnd0 ),
      .FSL3_S_EXISTS ( net_gnd0 ),
      .FSL3_M_CLK (  ),
      .FSL3_M_WRITE (  ),
      .FSL3_M_DATA (  ),
      .FSL3_M_CONTROL (  ),
      .FSL3_M_FULL ( net_gnd0 ),
      .FSL4_S_CLK (  ),
      .FSL4_S_READ (  ),
      .FSL4_S_DATA ( net_gnd32 ),
      .FSL4_S_CONTROL ( net_gnd0 ),
      .FSL4_S_EXISTS ( net_gnd0 ),
      .FSL4_M_CLK (  ),
      .FSL4_M_WRITE (  ),
      .FSL4_M_DATA (  ),
      .FSL4_M_CONTROL (  ),
      .FSL4_M_FULL ( net_gnd0 ),
      .FSL5_S_CLK (  ),
      .FSL5_S_READ (  ),
      .FSL5_S_DATA ( net_gnd32 ),
      .FSL5_S_CONTROL ( net_gnd0 ),
      .FSL5_S_EXISTS ( net_gnd0 ),
      .FSL5_M_CLK (  ),
      .FSL5_M_WRITE (  ),
      .FSL5_M_DATA (  ),
      .FSL5_M_CONTROL (  ),
      .FSL5_M_FULL ( net_gnd0 ),
      .FSL6_S_CLK (  ),
      .FSL6_S_READ (  ),
      .FSL6_S_DATA ( net_gnd32 ),
      .FSL6_S_CONTROL ( net_gnd0 ),
      .FSL6_S_EXISTS ( net_gnd0 ),
      .FSL6_M_CLK (  ),
      .FSL6_M_WRITE (  ),
      .FSL6_M_DATA (  ),
      .FSL6_M_CONTROL (  ),
      .FSL6_M_FULL ( net_gnd0 ),
      .FSL7_S_CLK (  ),
      .FSL7_S_READ (  ),
      .FSL7_S_DATA ( net_gnd32 ),
      .FSL7_S_CONTROL ( net_gnd0 ),
      .FSL7_S_EXISTS ( net_gnd0 ),
      .FSL7_M_CLK (  ),
      .FSL7_M_WRITE (  ),
      .FSL7_M_DATA (  ),
      .FSL7_M_CONTROL (  ),
      .FSL7_M_FULL ( net_gnd0 ),
      .FSL8_S_CLK (  ),
      .FSL8_S_READ (  ),
      .FSL8_S_DATA ( net_gnd32 ),
      .FSL8_S_CONTROL ( net_gnd0 ),
      .FSL8_S_EXISTS ( net_gnd0 ),
      .FSL8_M_CLK (  ),
      .FSL8_M_WRITE (  ),
      .FSL8_M_DATA (  ),
      .FSL8_M_CONTROL (  ),
      .FSL8_M_FULL ( net_gnd0 ),
      .FSL9_S_CLK (  ),
      .FSL9_S_READ (  ),
      .FSL9_S_DATA ( net_gnd32 ),
      .FSL9_S_CONTROL ( net_gnd0 ),
      .FSL9_S_EXISTS ( net_gnd0 ),
      .FSL9_M_CLK (  ),
      .FSL9_M_WRITE (  ),
      .FSL9_M_DATA (  ),
      .FSL9_M_CONTROL (  ),
      .FSL9_M_FULL ( net_gnd0 ),
      .FSL10_S_CLK (  ),
      .FSL10_S_READ (  ),
      .FSL10_S_DATA ( net_gnd32 ),
      .FSL10_S_CONTROL ( net_gnd0 ),
      .FSL10_S_EXISTS ( net_gnd0 ),
      .FSL10_M_CLK (  ),
      .FSL10_M_WRITE (  ),
      .FSL10_M_DATA (  ),
      .FSL10_M_CONTROL (  ),
      .FSL10_M_FULL ( net_gnd0 ),
      .FSL11_S_CLK (  ),
      .FSL11_S_READ (  ),
      .FSL11_S_DATA ( net_gnd32 ),
      .FSL11_S_CONTROL ( net_gnd0 ),
      .FSL11_S_EXISTS ( net_gnd0 ),
      .FSL11_M_CLK (  ),
      .FSL11_M_WRITE (  ),
      .FSL11_M_DATA (  ),
      .FSL11_M_CONTROL (  ),
      .FSL11_M_FULL ( net_gnd0 ),
      .FSL12_S_CLK (  ),
      .FSL12_S_READ (  ),
      .FSL12_S_DATA ( net_gnd32 ),
      .FSL12_S_CONTROL ( net_gnd0 ),
      .FSL12_S_EXISTS ( net_gnd0 ),
      .FSL12_M_CLK (  ),
      .FSL12_M_WRITE (  ),
      .FSL12_M_DATA (  ),
      .FSL12_M_CONTROL (  ),
      .FSL12_M_FULL ( net_gnd0 ),
      .FSL13_S_CLK (  ),
      .FSL13_S_READ (  ),
      .FSL13_S_DATA ( net_gnd32 ),
      .FSL13_S_CONTROL ( net_gnd0 ),
      .FSL13_S_EXISTS ( net_gnd0 ),
      .FSL13_M_CLK (  ),
      .FSL13_M_WRITE (  ),
      .FSL13_M_DATA (  ),
      .FSL13_M_CONTROL (  ),
      .FSL13_M_FULL ( net_gnd0 ),
      .FSL14_S_CLK (  ),
      .FSL14_S_READ (  ),
      .FSL14_S_DATA ( net_gnd32 ),
      .FSL14_S_CONTROL ( net_gnd0 ),
      .FSL14_S_EXISTS ( net_gnd0 ),
      .FSL14_M_CLK (  ),
      .FSL14_M_WRITE (  ),
      .FSL14_M_DATA (  ),
      .FSL14_M_CONTROL (  ),
      .FSL14_M_FULL ( net_gnd0 ),
      .FSL15_S_CLK (  ),
      .FSL15_S_READ (  ),
      .FSL15_S_DATA ( net_gnd32 ),
      .FSL15_S_CONTROL ( net_gnd0 ),
      .FSL15_S_EXISTS ( net_gnd0 ),
      .FSL15_M_CLK (  ),
      .FSL15_M_WRITE (  ),
      .FSL15_M_DATA (  ),
      .FSL15_M_CONTROL (  ),
      .FSL15_M_FULL ( net_gnd0 ),
      .M0_AXIS_TLAST (  ),
      .M0_AXIS_TDATA (  ),
      .M0_AXIS_TVALID (  ),
      .M0_AXIS_TREADY ( net_gnd0 ),
      .S0_AXIS_TLAST ( net_gnd0 ),
      .S0_AXIS_TDATA ( net_gnd32[0:31] ),
      .S0_AXIS_TVALID ( net_gnd0 ),
      .S0_AXIS_TREADY (  ),
      .M1_AXIS_TLAST (  ),
      .M1_AXIS_TDATA (  ),
      .M1_AXIS_TVALID (  ),
      .M1_AXIS_TREADY ( net_gnd0 ),
      .S1_AXIS_TLAST ( net_gnd0 ),
      .S1_AXIS_TDATA ( net_gnd32[0:31] ),
      .S1_AXIS_TVALID ( net_gnd0 ),
      .S1_AXIS_TREADY (  ),
      .M2_AXIS_TLAST (  ),
      .M2_AXIS_TDATA (  ),
      .M2_AXIS_TVALID (  ),
      .M2_AXIS_TREADY ( net_gnd0 ),
      .S2_AXIS_TLAST ( net_gnd0 ),
      .S2_AXIS_TDATA ( net_gnd32[0:31] ),
      .S2_AXIS_TVALID ( net_gnd0 ),
      .S2_AXIS_TREADY (  ),
      .M3_AXIS_TLAST (  ),
      .M3_AXIS_TDATA (  ),
      .M3_AXIS_TVALID (  ),
      .M3_AXIS_TREADY ( net_gnd0 ),
      .S3_AXIS_TLAST ( net_gnd0 ),
      .S3_AXIS_TDATA ( net_gnd32[0:31] ),
      .S3_AXIS_TVALID ( net_gnd0 ),
      .S3_AXIS_TREADY (  ),
      .M4_AXIS_TLAST (  ),
      .M4_AXIS_TDATA (  ),
      .M4_AXIS_TVALID (  ),
      .M4_AXIS_TREADY ( net_gnd0 ),
      .S4_AXIS_TLAST ( net_gnd0 ),
      .S4_AXIS_TDATA ( net_gnd32[0:31] ),
      .S4_AXIS_TVALID ( net_gnd0 ),
      .S4_AXIS_TREADY (  ),
      .M5_AXIS_TLAST (  ),
      .M5_AXIS_TDATA (  ),
      .M5_AXIS_TVALID (  ),
      .M5_AXIS_TREADY ( net_gnd0 ),
      .S5_AXIS_TLAST ( net_gnd0 ),
      .S5_AXIS_TDATA ( net_gnd32[0:31] ),
      .S5_AXIS_TVALID ( net_gnd0 ),
      .S5_AXIS_TREADY (  ),
      .M6_AXIS_TLAST (  ),
      .M6_AXIS_TDATA (  ),
      .M6_AXIS_TVALID (  ),
      .M6_AXIS_TREADY ( net_gnd0 ),
      .S6_AXIS_TLAST ( net_gnd0 ),
      .S6_AXIS_TDATA ( net_gnd32[0:31] ),
      .S6_AXIS_TVALID ( net_gnd0 ),
      .S6_AXIS_TREADY (  ),
      .M7_AXIS_TLAST (  ),
      .M7_AXIS_TDATA (  ),
      .M7_AXIS_TVALID (  ),
      .M7_AXIS_TREADY ( net_gnd0 ),
      .S7_AXIS_TLAST ( net_gnd0 ),
      .S7_AXIS_TDATA ( net_gnd32[0:31] ),
      .S7_AXIS_TVALID ( net_gnd0 ),
      .S7_AXIS_TREADY (  ),
      .M8_AXIS_TLAST (  ),
      .M8_AXIS_TDATA (  ),
      .M8_AXIS_TVALID (  ),
      .M8_AXIS_TREADY ( net_gnd0 ),
      .S8_AXIS_TLAST ( net_gnd0 ),
      .S8_AXIS_TDATA ( net_gnd32[0:31] ),
      .S8_AXIS_TVALID ( net_gnd0 ),
      .S8_AXIS_TREADY (  ),
      .M9_AXIS_TLAST (  ),
      .M9_AXIS_TDATA (  ),
      .M9_AXIS_TVALID (  ),
      .M9_AXIS_TREADY ( net_gnd0 ),
      .S9_AXIS_TLAST ( net_gnd0 ),
      .S9_AXIS_TDATA ( net_gnd32[0:31] ),
      .S9_AXIS_TVALID ( net_gnd0 ),
      .S9_AXIS_TREADY (  ),
      .M10_AXIS_TLAST (  ),
      .M10_AXIS_TDATA (  ),
      .M10_AXIS_TVALID (  ),
      .M10_AXIS_TREADY ( net_gnd0 ),
      .S10_AXIS_TLAST ( net_gnd0 ),
      .S10_AXIS_TDATA ( net_gnd32[0:31] ),
      .S10_AXIS_TVALID ( net_gnd0 ),
      .S10_AXIS_TREADY (  ),
      .M11_AXIS_TLAST (  ),
      .M11_AXIS_TDATA (  ),
      .M11_AXIS_TVALID (  ),
      .M11_AXIS_TREADY ( net_gnd0 ),
      .S11_AXIS_TLAST ( net_gnd0 ),
      .S11_AXIS_TDATA ( net_gnd32[0:31] ),
      .S11_AXIS_TVALID ( net_gnd0 ),
      .S11_AXIS_TREADY (  ),
      .M12_AXIS_TLAST (  ),
      .M12_AXIS_TDATA (  ),
      .M12_AXIS_TVALID (  ),
      .M12_AXIS_TREADY ( net_gnd0 ),
      .S12_AXIS_TLAST ( net_gnd0 ),
      .S12_AXIS_TDATA ( net_gnd32[0:31] ),
      .S12_AXIS_TVALID ( net_gnd0 ),
      .S12_AXIS_TREADY (  ),
      .M13_AXIS_TLAST (  ),
      .M13_AXIS_TDATA (  ),
      .M13_AXIS_TVALID (  ),
      .M13_AXIS_TREADY ( net_gnd0 ),
      .S13_AXIS_TLAST ( net_gnd0 ),
      .S13_AXIS_TDATA ( net_gnd32[0:31] ),
      .S13_AXIS_TVALID ( net_gnd0 ),
      .S13_AXIS_TREADY (  ),
      .M14_AXIS_TLAST (  ),
      .M14_AXIS_TDATA (  ),
      .M14_AXIS_TVALID (  ),
      .M14_AXIS_TREADY ( net_gnd0 ),
      .S14_AXIS_TLAST ( net_gnd0 ),
      .S14_AXIS_TDATA ( net_gnd32[0:31] ),
      .S14_AXIS_TVALID ( net_gnd0 ),
      .S14_AXIS_TREADY (  ),
      .M15_AXIS_TLAST (  ),
      .M15_AXIS_TDATA (  ),
      .M15_AXIS_TVALID (  ),
      .M15_AXIS_TREADY ( net_gnd0 ),
      .S15_AXIS_TLAST ( net_gnd0 ),
      .S15_AXIS_TDATA ( net_gnd32[0:31] ),
      .S15_AXIS_TVALID ( net_gnd0 ),
      .S15_AXIS_TREADY (  ),
      .ICACHE_FSL_IN_CLK (  ),
      .ICACHE_FSL_IN_READ (  ),
      .ICACHE_FSL_IN_DATA ( net_gnd32 ),
      .ICACHE_FSL_IN_CONTROL ( net_gnd0 ),
      .ICACHE_FSL_IN_EXISTS ( net_gnd0 ),
      .ICACHE_FSL_OUT_CLK (  ),
      .ICACHE_FSL_OUT_WRITE (  ),
      .ICACHE_FSL_OUT_DATA (  ),
      .ICACHE_FSL_OUT_CONTROL (  ),
      .ICACHE_FSL_OUT_FULL ( net_gnd0 ),
      .DCACHE_FSL_IN_CLK (  ),
      .DCACHE_FSL_IN_READ (  ),
      .DCACHE_FSL_IN_DATA ( net_gnd32 ),
      .DCACHE_FSL_IN_CONTROL ( net_gnd0 ),
      .DCACHE_FSL_IN_EXISTS ( net_gnd0 ),
      .DCACHE_FSL_OUT_CLK (  ),
      .DCACHE_FSL_OUT_WRITE (  ),
      .DCACHE_FSL_OUT_DATA (  ),
      .DCACHE_FSL_OUT_CONTROL (  ),
      .DCACHE_FSL_OUT_FULL ( net_gnd0 )
    );

  microblaze_mb_plb_wrapper
    mb_plb (
      .PLB_Clk ( clk_50_0000MHz ),
      .SYS_Rst ( sys_bus_reset[0] ),
      .PLB_Rst (  ),
      .SPLB_Rst ( mb_plb_SPLB_Rst ),
      .MPLB_Rst (  ),
      .PLB_dcrAck (  ),
      .PLB_dcrDBus (  ),
      .DCR_ABus ( net_gnd10 ),
      .DCR_DBus ( net_gnd32 ),
      .DCR_Read ( net_gnd0 ),
      .DCR_Write ( net_gnd0 ),
      .M_ABus ( mb_plb_M_ABus ),
      .M_UABus ( mb_plb_M_UABus ),
      .M_BE ( mb_plb_M_BE ),
      .M_RNW ( mb_plb_M_RNW ),
      .M_abort ( mb_plb_M_ABort ),
      .M_busLock ( mb_plb_M_busLock ),
      .M_TAttribute ( mb_plb_M_TAttribute ),
      .M_lockErr ( mb_plb_M_lockErr ),
      .M_MSize ( mb_plb_M_MSize ),
      .M_priority ( mb_plb_M_priority ),
      .M_rdBurst ( mb_plb_M_rdBurst ),
      .M_request ( mb_plb_M_request ),
      .M_size ( mb_plb_M_size ),
      .M_type ( mb_plb_M_type ),
      .M_wrBurst ( mb_plb_M_wrBurst ),
      .M_wrDBus ( mb_plb_M_wrDBus ),
      .Sl_addrAck ( mb_plb_Sl_addrAck ),
      .Sl_MRdErr ( mb_plb_Sl_MRdErr ),
      .Sl_MWrErr ( mb_plb_Sl_MWrErr ),
      .Sl_MBusy ( mb_plb_Sl_MBusy ),
      .Sl_rdBTerm ( mb_plb_Sl_rdBTerm ),
      .Sl_rdComp ( mb_plb_Sl_rdComp ),
      .Sl_rdDAck ( mb_plb_Sl_rdDAck ),
      .Sl_rdDBus ( mb_plb_Sl_rdDBus ),
      .Sl_rdWdAddr ( mb_plb_Sl_rdWdAddr ),
      .Sl_rearbitrate ( mb_plb_Sl_rearbitrate ),
      .Sl_SSize ( mb_plb_Sl_SSize ),
      .Sl_wait ( mb_plb_Sl_wait ),
      .Sl_wrBTerm ( mb_plb_Sl_wrBTerm ),
      .Sl_wrComp ( mb_plb_Sl_wrComp ),
      .Sl_wrDAck ( mb_plb_Sl_wrDAck ),
      .Sl_MIRQ ( mb_plb_Sl_MIRQ ),
      .PLB_MIRQ ( mb_plb_PLB_MIRQ ),
      .PLB_ABus ( mb_plb_PLB_ABus ),
      .PLB_UABus ( mb_plb_PLB_UABus ),
      .PLB_BE ( mb_plb_PLB_BE ),
      .PLB_MAddrAck ( mb_plb_PLB_MAddrAck ),
      .PLB_MTimeout ( mb_plb_PLB_MTimeout ),
      .PLB_MBusy ( mb_plb_PLB_MBusy ),
      .PLB_MRdErr ( mb_plb_PLB_MRdErr ),
      .PLB_MWrErr ( mb_plb_PLB_MWrErr ),
      .PLB_MRdBTerm ( mb_plb_PLB_MRdBTerm ),
      .PLB_MRdDAck ( mb_plb_PLB_MRdDAck ),
      .PLB_MRdDBus ( mb_plb_PLB_MRdDBus ),
      .PLB_MRdWdAddr ( mb_plb_PLB_MRdWdAddr ),
      .PLB_MRearbitrate ( mb_plb_PLB_MRearbitrate ),
      .PLB_MWrBTerm ( mb_plb_PLB_MWrBTerm ),
      .PLB_MWrDAck ( mb_plb_PLB_MWrDAck ),
      .PLB_MSSize ( mb_plb_PLB_MSSize ),
      .PLB_PAValid ( mb_plb_PLB_PAValid ),
      .PLB_RNW ( mb_plb_PLB_RNW ),
      .PLB_SAValid ( mb_plb_PLB_SAValid ),
      .PLB_abort ( mb_plb_PLB_abort ),
      .PLB_busLock ( mb_plb_PLB_busLock ),
      .PLB_TAttribute ( mb_plb_PLB_TAttribute ),
      .PLB_lockErr ( mb_plb_PLB_lockErr ),
      .PLB_masterID ( mb_plb_PLB_masterID[0:0] ),
      .PLB_MSize ( mb_plb_PLB_MSize ),
      .PLB_rdPendPri ( mb_plb_PLB_rdPendPri ),
      .PLB_wrPendPri ( mb_plb_PLB_wrPendPri ),
      .PLB_rdPendReq ( mb_plb_PLB_rdPendReq ),
      .PLB_wrPendReq ( mb_plb_PLB_wrPendReq ),
      .PLB_rdBurst ( mb_plb_PLB_rdBurst ),
      .PLB_rdPrim ( mb_plb_PLB_rdPrim ),
      .PLB_reqPri ( mb_plb_PLB_reqPri ),
      .PLB_size ( mb_plb_PLB_size ),
      .PLB_type ( mb_plb_PLB_type ),
      .PLB_wrBurst ( mb_plb_PLB_wrBurst ),
      .PLB_wrDBus ( mb_plb_PLB_wrDBus ),
      .PLB_wrPrim ( mb_plb_PLB_wrPrim ),
      .PLB_SaddrAck (  ),
      .PLB_SMRdErr (  ),
      .PLB_SMWrErr (  ),
      .PLB_SMBusy (  ),
      .PLB_SrdBTerm (  ),
      .PLB_SrdComp (  ),
      .PLB_SrdDAck (  ),
      .PLB_SrdDBus (  ),
      .PLB_SrdWdAddr (  ),
      .PLB_Srearbitrate (  ),
      .PLB_Sssize (  ),
      .PLB_Swait (  ),
      .PLB_SwrBTerm (  ),
      .PLB_SwrComp (  ),
      .PLB_SwrDAck (  ),
      .Bus_Error_Det (  )
    );

  microblaze_ilmb_wrapper
    ilmb (
      .LMB_Clk ( clk_50_0000MHz ),
      .SYS_Rst ( sys_bus_reset[0] ),
      .LMB_Rst ( ilmb_LMB_Rst ),
      .M_ABus ( ilmb_M_ABus ),
      .M_ReadStrobe ( ilmb_M_ReadStrobe ),
      .M_WriteStrobe ( net_gnd0 ),
      .M_AddrStrobe ( ilmb_M_AddrStrobe ),
      .M_DBus ( net_gnd32 ),
      .M_BE ( net_gnd4 ),
      .Sl_DBus ( ilmb_Sl_DBus ),
      .Sl_Ready ( ilmb_Sl_Ready[0:0] ),
      .Sl_Wait ( ilmb_Sl_Wait[0:0] ),
      .Sl_UE ( ilmb_Sl_UE[0:0] ),
      .Sl_CE ( ilmb_Sl_CE[0:0] ),
      .LMB_ABus ( ilmb_LMB_ABus ),
      .LMB_ReadStrobe ( ilmb_LMB_ReadStrobe ),
      .LMB_WriteStrobe ( ilmb_LMB_WriteStrobe ),
      .LMB_AddrStrobe ( ilmb_LMB_AddrStrobe ),
      .LMB_ReadDBus ( ilmb_LMB_ReadDBus ),
      .LMB_WriteDBus ( ilmb_LMB_WriteDBus ),
      .LMB_Ready ( ilmb_LMB_Ready ),
      .LMB_Wait ( ilmb_LMB_Wait ),
      .LMB_UE ( ilmb_LMB_UE ),
      .LMB_CE ( ilmb_LMB_CE ),
      .LMB_BE ( ilmb_LMB_BE )
    );

  microblaze_dlmb_wrapper
    dlmb (
      .LMB_Clk ( clk_50_0000MHz ),
      .SYS_Rst ( sys_bus_reset[0] ),
      .LMB_Rst ( dlmb_LMB_Rst ),
      .M_ABus ( dlmb_M_ABus ),
      .M_ReadStrobe ( dlmb_M_ReadStrobe ),
      .M_WriteStrobe ( dlmb_M_WriteStrobe ),
      .M_AddrStrobe ( dlmb_M_AddrStrobe ),
      .M_DBus ( dlmb_M_DBus ),
      .M_BE ( dlmb_M_BE ),
      .Sl_DBus ( dlmb_Sl_DBus ),
      .Sl_Ready ( dlmb_Sl_Ready[0:0] ),
      .Sl_Wait ( dlmb_Sl_Wait[0:0] ),
      .Sl_UE ( dlmb_Sl_UE[0:0] ),
      .Sl_CE ( dlmb_Sl_CE[0:0] ),
      .LMB_ABus ( dlmb_LMB_ABus ),
      .LMB_ReadStrobe ( dlmb_LMB_ReadStrobe ),
      .LMB_WriteStrobe ( dlmb_LMB_WriteStrobe ),
      .LMB_AddrStrobe ( dlmb_LMB_AddrStrobe ),
      .LMB_ReadDBus ( dlmb_LMB_ReadDBus ),
      .LMB_WriteDBus ( dlmb_LMB_WriteDBus ),
      .LMB_Ready ( dlmb_LMB_Ready ),
      .LMB_Wait ( dlmb_LMB_Wait ),
      .LMB_UE ( dlmb_LMB_UE ),
      .LMB_CE ( dlmb_LMB_CE ),
      .LMB_BE ( dlmb_LMB_BE )
    );

  microblaze_dlmb_cntlr_wrapper
    dlmb_cntlr (
      .LMB_Clk ( clk_50_0000MHz ),
      .LMB_Rst ( dlmb_LMB_Rst ),
      .LMB_ABus ( dlmb_LMB_ABus ),
      .LMB_WriteDBus ( dlmb_LMB_WriteDBus ),
      .LMB_AddrStrobe ( dlmb_LMB_AddrStrobe ),
      .LMB_ReadStrobe ( dlmb_LMB_ReadStrobe ),
      .LMB_WriteStrobe ( dlmb_LMB_WriteStrobe ),
      .LMB_BE ( dlmb_LMB_BE ),
      .Sl_DBus ( dlmb_Sl_DBus ),
      .Sl_Ready ( dlmb_Sl_Ready[0] ),
      .Sl_Wait ( dlmb_Sl_Wait[0] ),
      .Sl_UE ( dlmb_Sl_UE[0] ),
      .Sl_CE ( dlmb_Sl_CE[0] ),
      .LMB1_ABus ( net_gnd32 ),
      .LMB1_WriteDBus ( net_gnd32 ),
      .LMB1_AddrStrobe ( net_gnd0 ),
      .LMB1_ReadStrobe ( net_gnd0 ),
      .LMB1_WriteStrobe ( net_gnd0 ),
      .LMB1_BE ( net_gnd4 ),
      .Sl1_DBus (  ),
      .Sl1_Ready (  ),
      .Sl1_Wait (  ),
      .Sl1_UE (  ),
      .Sl1_CE (  ),
      .LMB2_ABus ( net_gnd32 ),
      .LMB2_WriteDBus ( net_gnd32 ),
      .LMB2_AddrStrobe ( net_gnd0 ),
      .LMB2_ReadStrobe ( net_gnd0 ),
      .LMB2_WriteStrobe ( net_gnd0 ),
      .LMB2_BE ( net_gnd4 ),
      .Sl2_DBus (  ),
      .Sl2_Ready (  ),
      .Sl2_Wait (  ),
      .Sl2_UE (  ),
      .Sl2_CE (  ),
      .LMB3_ABus ( net_gnd32 ),
      .LMB3_WriteDBus ( net_gnd32 ),
      .LMB3_AddrStrobe ( net_gnd0 ),
      .LMB3_ReadStrobe ( net_gnd0 ),
      .LMB3_WriteStrobe ( net_gnd0 ),
      .LMB3_BE ( net_gnd4 ),
      .Sl3_DBus (  ),
      .Sl3_Ready (  ),
      .Sl3_Wait (  ),
      .Sl3_UE (  ),
      .Sl3_CE (  ),
      .BRAM_Rst_A ( dlmb_port_BRAM_Rst ),
      .BRAM_Clk_A ( dlmb_port_BRAM_Clk ),
      .BRAM_EN_A ( dlmb_port_BRAM_EN ),
      .BRAM_WEN_A ( dlmb_port_BRAM_WEN ),
      .BRAM_Addr_A ( dlmb_port_BRAM_Addr ),
      .BRAM_Din_A ( dlmb_port_BRAM_Din ),
      .BRAM_Dout_A ( dlmb_port_BRAM_Dout ),
      .Interrupt (  ),
      .UE (  ),
      .CE (  ),
      .SPLB_CTRL_PLB_ABus ( net_gnd32 ),
      .SPLB_CTRL_PLB_PAValid ( net_gnd0 ),
      .SPLB_CTRL_PLB_masterID ( net_gnd1[0:0] ),
      .SPLB_CTRL_PLB_RNW ( net_gnd0 ),
      .SPLB_CTRL_PLB_BE ( net_gnd4 ),
      .SPLB_CTRL_PLB_size ( net_gnd4 ),
      .SPLB_CTRL_PLB_type ( net_gnd3[2:0] ),
      .SPLB_CTRL_PLB_wrDBus ( net_gnd32 ),
      .SPLB_CTRL_Sl_addrAck (  ),
      .SPLB_CTRL_Sl_SSize (  ),
      .SPLB_CTRL_Sl_wait (  ),
      .SPLB_CTRL_Sl_rearbitrate (  ),
      .SPLB_CTRL_Sl_wrDAck (  ),
      .SPLB_CTRL_Sl_wrComp (  ),
      .SPLB_CTRL_Sl_rdDBus (  ),
      .SPLB_CTRL_Sl_rdDAck (  ),
      .SPLB_CTRL_Sl_rdComp (  ),
      .SPLB_CTRL_Sl_MBusy (  ),
      .SPLB_CTRL_Sl_MWrErr (  ),
      .SPLB_CTRL_Sl_MRdErr (  ),
      .SPLB_CTRL_PLB_UABus ( net_gnd32 ),
      .SPLB_CTRL_PLB_SAValid ( net_gnd0 ),
      .SPLB_CTRL_PLB_rdPrim ( net_gnd0 ),
      .SPLB_CTRL_PLB_wrPrim ( net_gnd0 ),
      .SPLB_CTRL_PLB_abort ( net_gnd0 ),
      .SPLB_CTRL_PLB_busLock ( net_gnd0 ),
      .SPLB_CTRL_PLB_MSize ( net_gnd2 ),
      .SPLB_CTRL_PLB_lockErr ( net_gnd0 ),
      .SPLB_CTRL_PLB_wrBurst ( net_gnd0 ),
      .SPLB_CTRL_PLB_rdBurst ( net_gnd0 ),
      .SPLB_CTRL_PLB_wrPendReq ( net_gnd0 ),
      .SPLB_CTRL_PLB_rdPendReq ( net_gnd0 ),
      .SPLB_CTRL_PLB_wrPendPri ( net_gnd2 ),
      .SPLB_CTRL_PLB_rdPendPri ( net_gnd2 ),
      .SPLB_CTRL_PLB_reqPri ( net_gnd2 ),
      .SPLB_CTRL_PLB_TAttribute ( net_gnd16 ),
      .SPLB_CTRL_Sl_wrBTerm (  ),
      .SPLB_CTRL_Sl_rdWdAddr (  ),
      .SPLB_CTRL_Sl_rdBTerm (  ),
      .SPLB_CTRL_Sl_MIRQ (  ),
      .S_AXI_CTRL_ACLK ( net_vcc0 ),
      .S_AXI_CTRL_ARESETN ( net_gnd0 ),
      .S_AXI_CTRL_AWADDR ( net_gnd32[0:31] ),
      .S_AXI_CTRL_AWVALID ( net_gnd0 ),
      .S_AXI_CTRL_AWREADY (  ),
      .S_AXI_CTRL_WDATA ( net_gnd32[0:31] ),
      .S_AXI_CTRL_WSTRB ( net_gnd4[0:3] ),
      .S_AXI_CTRL_WVALID ( net_gnd0 ),
      .S_AXI_CTRL_WREADY (  ),
      .S_AXI_CTRL_BRESP (  ),
      .S_AXI_CTRL_BVALID (  ),
      .S_AXI_CTRL_BREADY ( net_gnd0 ),
      .S_AXI_CTRL_ARADDR ( net_gnd32[0:31] ),
      .S_AXI_CTRL_ARVALID ( net_gnd0 ),
      .S_AXI_CTRL_ARREADY (  ),
      .S_AXI_CTRL_RDATA (  ),
      .S_AXI_CTRL_RRESP (  ),
      .S_AXI_CTRL_RVALID (  ),
      .S_AXI_CTRL_RREADY ( net_gnd0 )
    );

  microblaze_ilmb_cntlr_wrapper
    ilmb_cntlr (
      .LMB_Clk ( clk_50_0000MHz ),
      .LMB_Rst ( ilmb_LMB_Rst ),
      .LMB_ABus ( ilmb_LMB_ABus ),
      .LMB_WriteDBus ( ilmb_LMB_WriteDBus ),
      .LMB_AddrStrobe ( ilmb_LMB_AddrStrobe ),
      .LMB_ReadStrobe ( ilmb_LMB_ReadStrobe ),
      .LMB_WriteStrobe ( ilmb_LMB_WriteStrobe ),
      .LMB_BE ( ilmb_LMB_BE ),
      .Sl_DBus ( ilmb_Sl_DBus ),
      .Sl_Ready ( ilmb_Sl_Ready[0] ),
      .Sl_Wait ( ilmb_Sl_Wait[0] ),
      .Sl_UE ( ilmb_Sl_UE[0] ),
      .Sl_CE ( ilmb_Sl_CE[0] ),
      .LMB1_ABus ( net_gnd32 ),
      .LMB1_WriteDBus ( net_gnd32 ),
      .LMB1_AddrStrobe ( net_gnd0 ),
      .LMB1_ReadStrobe ( net_gnd0 ),
      .LMB1_WriteStrobe ( net_gnd0 ),
      .LMB1_BE ( net_gnd4 ),
      .Sl1_DBus (  ),
      .Sl1_Ready (  ),
      .Sl1_Wait (  ),
      .Sl1_UE (  ),
      .Sl1_CE (  ),
      .LMB2_ABus ( net_gnd32 ),
      .LMB2_WriteDBus ( net_gnd32 ),
      .LMB2_AddrStrobe ( net_gnd0 ),
      .LMB2_ReadStrobe ( net_gnd0 ),
      .LMB2_WriteStrobe ( net_gnd0 ),
      .LMB2_BE ( net_gnd4 ),
      .Sl2_DBus (  ),
      .Sl2_Ready (  ),
      .Sl2_Wait (  ),
      .Sl2_UE (  ),
      .Sl2_CE (  ),
      .LMB3_ABus ( net_gnd32 ),
      .LMB3_WriteDBus ( net_gnd32 ),
      .LMB3_AddrStrobe ( net_gnd0 ),
      .LMB3_ReadStrobe ( net_gnd0 ),
      .LMB3_WriteStrobe ( net_gnd0 ),
      .LMB3_BE ( net_gnd4 ),
      .Sl3_DBus (  ),
      .Sl3_Ready (  ),
      .Sl3_Wait (  ),
      .Sl3_UE (  ),
      .Sl3_CE (  ),
      .BRAM_Rst_A ( ilmb_cntlr_BRAM_PORT_BRAM_Rst ),
      .BRAM_Clk_A ( ilmb_cntlr_BRAM_PORT_BRAM_Clk ),
      .BRAM_EN_A ( ilmb_cntlr_BRAM_PORT_BRAM_EN ),
      .BRAM_WEN_A ( ilmb_cntlr_BRAM_PORT_BRAM_WEN ),
      .BRAM_Addr_A ( ilmb_cntlr_BRAM_PORT_BRAM_Addr ),
      .BRAM_Din_A ( ilmb_cntlr_BRAM_PORT_BRAM_Din ),
      .BRAM_Dout_A ( ilmb_cntlr_BRAM_PORT_BRAM_Dout ),
      .Interrupt (  ),
      .UE (  ),
      .CE (  ),
      .SPLB_CTRL_PLB_ABus ( net_gnd32 ),
      .SPLB_CTRL_PLB_PAValid ( net_gnd0 ),
      .SPLB_CTRL_PLB_masterID ( net_gnd1[0:0] ),
      .SPLB_CTRL_PLB_RNW ( net_gnd0 ),
      .SPLB_CTRL_PLB_BE ( net_gnd4 ),
      .SPLB_CTRL_PLB_size ( net_gnd4 ),
      .SPLB_CTRL_PLB_type ( net_gnd3[2:0] ),
      .SPLB_CTRL_PLB_wrDBus ( net_gnd32 ),
      .SPLB_CTRL_Sl_addrAck (  ),
      .SPLB_CTRL_Sl_SSize (  ),
      .SPLB_CTRL_Sl_wait (  ),
      .SPLB_CTRL_Sl_rearbitrate (  ),
      .SPLB_CTRL_Sl_wrDAck (  ),
      .SPLB_CTRL_Sl_wrComp (  ),
      .SPLB_CTRL_Sl_rdDBus (  ),
      .SPLB_CTRL_Sl_rdDAck (  ),
      .SPLB_CTRL_Sl_rdComp (  ),
      .SPLB_CTRL_Sl_MBusy (  ),
      .SPLB_CTRL_Sl_MWrErr (  ),
      .SPLB_CTRL_Sl_MRdErr (  ),
      .SPLB_CTRL_PLB_UABus ( net_gnd32 ),
      .SPLB_CTRL_PLB_SAValid ( net_gnd0 ),
      .SPLB_CTRL_PLB_rdPrim ( net_gnd0 ),
      .SPLB_CTRL_PLB_wrPrim ( net_gnd0 ),
      .SPLB_CTRL_PLB_abort ( net_gnd0 ),
      .SPLB_CTRL_PLB_busLock ( net_gnd0 ),
      .SPLB_CTRL_PLB_MSize ( net_gnd2 ),
      .SPLB_CTRL_PLB_lockErr ( net_gnd0 ),
      .SPLB_CTRL_PLB_wrBurst ( net_gnd0 ),
      .SPLB_CTRL_PLB_rdBurst ( net_gnd0 ),
      .SPLB_CTRL_PLB_wrPendReq ( net_gnd0 ),
      .SPLB_CTRL_PLB_rdPendReq ( net_gnd0 ),
      .SPLB_CTRL_PLB_wrPendPri ( net_gnd2 ),
      .SPLB_CTRL_PLB_rdPendPri ( net_gnd2 ),
      .SPLB_CTRL_PLB_reqPri ( net_gnd2 ),
      .SPLB_CTRL_PLB_TAttribute ( net_gnd16 ),
      .SPLB_CTRL_Sl_wrBTerm (  ),
      .SPLB_CTRL_Sl_rdWdAddr (  ),
      .SPLB_CTRL_Sl_rdBTerm (  ),
      .SPLB_CTRL_Sl_MIRQ (  ),
      .S_AXI_CTRL_ACLK ( net_vcc0 ),
      .S_AXI_CTRL_ARESETN ( net_gnd0 ),
      .S_AXI_CTRL_AWADDR ( net_gnd32[0:31] ),
      .S_AXI_CTRL_AWVALID ( net_gnd0 ),
      .S_AXI_CTRL_AWREADY (  ),
      .S_AXI_CTRL_WDATA ( net_gnd32[0:31] ),
      .S_AXI_CTRL_WSTRB ( net_gnd4[0:3] ),
      .S_AXI_CTRL_WVALID ( net_gnd0 ),
      .S_AXI_CTRL_WREADY (  ),
      .S_AXI_CTRL_BRESP (  ),
      .S_AXI_CTRL_BVALID (  ),
      .S_AXI_CTRL_BREADY ( net_gnd0 ),
      .S_AXI_CTRL_ARADDR ( net_gnd32[0:31] ),
      .S_AXI_CTRL_ARVALID ( net_gnd0 ),
      .S_AXI_CTRL_ARREADY (  ),
      .S_AXI_CTRL_RDATA (  ),
      .S_AXI_CTRL_RRESP (  ),
      .S_AXI_CTRL_RVALID (  ),
      .S_AXI_CTRL_RREADY ( net_gnd0 )
    );

  microblaze_lmb_bram_wrapper
    lmb_bram (
      .BRAM_Rst_A ( dlmb_port_BRAM_Rst ),
      .BRAM_Clk_A ( dlmb_port_BRAM_Clk ),
      .BRAM_EN_A ( dlmb_port_BRAM_EN ),
      .BRAM_WEN_A ( dlmb_port_BRAM_WEN ),
      .BRAM_Addr_A ( dlmb_port_BRAM_Addr ),
      .BRAM_Din_A ( dlmb_port_BRAM_Din ),
      .BRAM_Dout_A ( dlmb_port_BRAM_Dout ),
      .BRAM_Rst_B ( ilmb_cntlr_BRAM_PORT_BRAM_Rst ),
      .BRAM_Clk_B ( ilmb_cntlr_BRAM_PORT_BRAM_Clk ),
      .BRAM_EN_B ( ilmb_cntlr_BRAM_PORT_BRAM_EN ),
      .BRAM_WEN_B ( ilmb_cntlr_BRAM_PORT_BRAM_WEN ),
      .BRAM_Addr_B ( ilmb_cntlr_BRAM_PORT_BRAM_Addr ),
      .BRAM_Din_B ( ilmb_cntlr_BRAM_PORT_BRAM_Din ),
      .BRAM_Dout_B ( ilmb_cntlr_BRAM_PORT_BRAM_Dout )
    );

  microblaze_rs232_wrapper
    RS232 (
      .SPLB_Clk ( clk_50_0000MHz ),
      .SPLB_Rst ( mb_plb_SPLB_Rst[0] ),
      .PLB_ABus ( mb_plb_PLB_ABus ),
      .PLB_PAValid ( mb_plb_PLB_PAValid ),
      .PLB_masterID ( mb_plb_PLB_masterID[0:0] ),
      .PLB_RNW ( mb_plb_PLB_RNW ),
      .PLB_BE ( mb_plb_PLB_BE ),
      .PLB_size ( mb_plb_PLB_size ),
      .PLB_type ( mb_plb_PLB_type ),
      .PLB_wrDBus ( mb_plb_PLB_wrDBus ),
      .PLB_UABus ( mb_plb_PLB_UABus ),
      .PLB_SAValid ( mb_plb_PLB_SAValid ),
      .PLB_rdPrim ( mb_plb_PLB_rdPrim[0] ),
      .PLB_wrPrim ( mb_plb_PLB_wrPrim[0] ),
      .PLB_abort ( mb_plb_PLB_abort ),
      .PLB_busLock ( mb_plb_PLB_busLock ),
      .PLB_MSize ( mb_plb_PLB_MSize ),
      .PLB_lockErr ( mb_plb_PLB_lockErr ),
      .PLB_wrBurst ( mb_plb_PLB_wrBurst ),
      .PLB_rdBurst ( mb_plb_PLB_rdBurst ),
      .PLB_wrPendReq ( mb_plb_PLB_wrPendReq ),
      .PLB_rdPendReq ( mb_plb_PLB_rdPendReq ),
      .PLB_wrPendPri ( mb_plb_PLB_wrPendPri ),
      .PLB_rdPendPri ( mb_plb_PLB_rdPendPri ),
      .PLB_reqPri ( mb_plb_PLB_reqPri ),
      .PLB_TAttribute ( mb_plb_PLB_TAttribute ),
      .Sl_addrAck ( mb_plb_Sl_addrAck[0] ),
      .Sl_SSize ( mb_plb_Sl_SSize[0:1] ),
      .Sl_wait ( mb_plb_Sl_wait[0] ),
      .Sl_rearbitrate ( mb_plb_Sl_rearbitrate[0] ),
      .Sl_wrDAck ( mb_plb_Sl_wrDAck[0] ),
      .Sl_wrComp ( mb_plb_Sl_wrComp[0] ),
      .Sl_rdDBus ( mb_plb_Sl_rdDBus[0:31] ),
      .Sl_rdDAck ( mb_plb_Sl_rdDAck[0] ),
      .Sl_rdComp ( mb_plb_Sl_rdComp[0] ),
      .Sl_MBusy ( mb_plb_Sl_MBusy[0:1] ),
      .Sl_MWrErr ( mb_plb_Sl_MWrErr[0:1] ),
      .Sl_MRdErr ( mb_plb_Sl_MRdErr[0:1] ),
      .Sl_wrBTerm ( mb_plb_Sl_wrBTerm[0] ),
      .Sl_rdWdAddr ( mb_plb_Sl_rdWdAddr[0:3] ),
      .Sl_rdBTerm ( mb_plb_Sl_rdBTerm[0] ),
      .Sl_MIRQ ( mb_plb_Sl_MIRQ[0:1] ),
      .RX ( fpga_0_RS232_RX_pin ),
      .TX ( fpga_0_RS232_TX_pin ),
      .Interrupt ( RS232_Interrupt[0] )
    );

  microblaze_clock_generator_0_wrapper
    clock_generator_0 (
      .CLKIN ( CLK_S ),
      .CLKOUT0 ( clk_50_0000MHz ),
      .CLKOUT1 (  ),
      .CLKOUT2 (  ),
      .CLKOUT3 (  ),
      .CLKOUT4 (  ),
      .CLKOUT5 (  ),
      .CLKOUT6 (  ),
      .CLKOUT7 (  ),
      .CLKOUT8 (  ),
      .CLKOUT9 (  ),
      .CLKOUT10 (  ),
      .CLKOUT11 (  ),
      .CLKOUT12 (  ),
      .CLKOUT13 (  ),
      .CLKOUT14 (  ),
      .CLKOUT15 (  ),
      .CLKFBIN ( net_gnd0 ),
      .CLKFBOUT (  ),
      .PSCLK ( net_gnd0 ),
      .PSEN ( net_gnd0 ),
      .PSINCDEC ( net_gnd0 ),
      .PSDONE (  ),
      .RST ( sys_rst_s ),
      .LOCKED ( Dcm_all_locked )
    );

  microblaze_mdm_0_wrapper
    mdm_0 (
      .Interrupt (  ),
      .Debug_SYS_Rst ( Debug_SYS_Rst ),
      .Ext_BRK ( Ext_BRK ),
      .Ext_NM_BRK ( Ext_NM_BRK ),
      .S_AXI_ACLK ( net_gnd0 ),
      .S_AXI_ARESETN ( net_gnd0 ),
      .S_AXI_AWADDR ( net_gnd32[0:31] ),
      .S_AXI_AWVALID ( net_gnd0 ),
      .S_AXI_AWREADY (  ),
      .S_AXI_WDATA ( net_gnd32[0:31] ),
      .S_AXI_WSTRB ( net_gnd4[0:3] ),
      .S_AXI_WVALID ( net_gnd0 ),
      .S_AXI_WREADY (  ),
      .S_AXI_BRESP (  ),
      .S_AXI_BVALID (  ),
      .S_AXI_BREADY ( net_gnd0 ),
      .S_AXI_ARADDR ( net_gnd32[0:31] ),
      .S_AXI_ARVALID ( net_gnd0 ),
      .S_AXI_ARREADY (  ),
      .S_AXI_RDATA (  ),
      .S_AXI_RRESP (  ),
      .S_AXI_RVALID (  ),
      .S_AXI_RREADY ( net_gnd0 ),
      .SPLB_Clk ( clk_50_0000MHz ),
      .SPLB_Rst ( mb_plb_SPLB_Rst[1] ),
      .PLB_ABus ( mb_plb_PLB_ABus ),
      .PLB_UABus ( mb_plb_PLB_UABus ),
      .PLB_PAValid ( mb_plb_PLB_PAValid ),
      .PLB_SAValid ( mb_plb_PLB_SAValid ),
      .PLB_rdPrim ( mb_plb_PLB_rdPrim[1] ),
      .PLB_wrPrim ( mb_plb_PLB_wrPrim[1] ),
      .PLB_masterID ( mb_plb_PLB_masterID[0:0] ),
      .PLB_abort ( mb_plb_PLB_abort ),
      .PLB_busLock ( mb_plb_PLB_busLock ),
      .PLB_RNW ( mb_plb_PLB_RNW ),
      .PLB_BE ( mb_plb_PLB_BE ),
      .PLB_MSize ( mb_plb_PLB_MSize ),
      .PLB_size ( mb_plb_PLB_size ),
      .PLB_type ( mb_plb_PLB_type ),
      .PLB_lockErr ( mb_plb_PLB_lockErr ),
      .PLB_wrDBus ( mb_plb_PLB_wrDBus ),
      .PLB_wrBurst ( mb_plb_PLB_wrBurst ),
      .PLB_rdBurst ( mb_plb_PLB_rdBurst ),
      .PLB_wrPendReq ( mb_plb_PLB_wrPendReq ),
      .PLB_rdPendReq ( mb_plb_PLB_rdPendReq ),
      .PLB_wrPendPri ( mb_plb_PLB_wrPendPri ),
      .PLB_rdPendPri ( mb_plb_PLB_rdPendPri ),
      .PLB_reqPri ( mb_plb_PLB_reqPri ),
      .PLB_TAttribute ( mb_plb_PLB_TAttribute ),
      .Sl_addrAck ( mb_plb_Sl_addrAck[1] ),
      .Sl_SSize ( mb_plb_Sl_SSize[2:3] ),
      .Sl_wait ( mb_plb_Sl_wait[1] ),
      .Sl_rearbitrate ( mb_plb_Sl_rearbitrate[1] ),
      .Sl_wrDAck ( mb_plb_Sl_wrDAck[1] ),
      .Sl_wrComp ( mb_plb_Sl_wrComp[1] ),
      .Sl_wrBTerm ( mb_plb_Sl_wrBTerm[1] ),
      .Sl_rdDBus ( mb_plb_Sl_rdDBus[32:63] ),
      .Sl_rdWdAddr ( mb_plb_Sl_rdWdAddr[4:7] ),
      .Sl_rdDAck ( mb_plb_Sl_rdDAck[1] ),
      .Sl_rdComp ( mb_plb_Sl_rdComp[1] ),
      .Sl_rdBTerm ( mb_plb_Sl_rdBTerm[1] ),
      .Sl_MBusy ( mb_plb_Sl_MBusy[2:3] ),
      .Sl_MWrErr ( mb_plb_Sl_MWrErr[2:3] ),
      .Sl_MRdErr ( mb_plb_Sl_MRdErr[2:3] ),
      .Sl_MIRQ ( mb_plb_Sl_MIRQ[2:3] ),
      .Dbg_Clk_0 ( microblaze_0_mdm_bus_Dbg_Clk ),
      .Dbg_TDI_0 ( microblaze_0_mdm_bus_Dbg_TDI ),
      .Dbg_TDO_0 ( microblaze_0_mdm_bus_Dbg_TDO ),
      .Dbg_Reg_En_0 ( microblaze_0_mdm_bus_Dbg_Reg_En ),
      .Dbg_Capture_0 ( microblaze_0_mdm_bus_Dbg_Capture ),
      .Dbg_Shift_0 ( microblaze_0_mdm_bus_Dbg_Shift ),
      .Dbg_Update_0 ( microblaze_0_mdm_bus_Dbg_Update ),
      .Dbg_Rst_0 ( microblaze_0_mdm_bus_Debug_Rst ),
      .Dbg_Clk_1 (  ),
      .Dbg_TDI_1 (  ),
      .Dbg_TDO_1 ( net_gnd0 ),
      .Dbg_Reg_En_1 (  ),
      .Dbg_Capture_1 (  ),
      .Dbg_Shift_1 (  ),
      .Dbg_Update_1 (  ),
      .Dbg_Rst_1 (  ),
      .Dbg_Clk_2 (  ),
      .Dbg_TDI_2 (  ),
      .Dbg_TDO_2 ( net_gnd0 ),
      .Dbg_Reg_En_2 (  ),
      .Dbg_Capture_2 (  ),
      .Dbg_Shift_2 (  ),
      .Dbg_Update_2 (  ),
      .Dbg_Rst_2 (  ),
      .Dbg_Clk_3 (  ),
      .Dbg_TDI_3 (  ),
      .Dbg_TDO_3 ( net_gnd0 ),
      .Dbg_Reg_En_3 (  ),
      .Dbg_Capture_3 (  ),
      .Dbg_Shift_3 (  ),
      .Dbg_Update_3 (  ),
      .Dbg_Rst_3 (  ),
      .Dbg_Clk_4 (  ),
      .Dbg_TDI_4 (  ),
      .Dbg_TDO_4 ( net_gnd0 ),
      .Dbg_Reg_En_4 (  ),
      .Dbg_Capture_4 (  ),
      .Dbg_Shift_4 (  ),
      .Dbg_Update_4 (  ),
      .Dbg_Rst_4 (  ),
      .Dbg_Clk_5 (  ),
      .Dbg_TDI_5 (  ),
      .Dbg_TDO_5 ( net_gnd0 ),
      .Dbg_Reg_En_5 (  ),
      .Dbg_Capture_5 (  ),
      .Dbg_Shift_5 (  ),
      .Dbg_Update_5 (  ),
      .Dbg_Rst_5 (  ),
      .Dbg_Clk_6 (  ),
      .Dbg_TDI_6 (  ),
      .Dbg_TDO_6 ( net_gnd0 ),
      .Dbg_Reg_En_6 (  ),
      .Dbg_Capture_6 (  ),
      .Dbg_Shift_6 (  ),
      .Dbg_Update_6 (  ),
      .Dbg_Rst_6 (  ),
      .Dbg_Clk_7 (  ),
      .Dbg_TDI_7 (  ),
      .Dbg_TDO_7 ( net_gnd0 ),
      .Dbg_Reg_En_7 (  ),
      .Dbg_Capture_7 (  ),
      .Dbg_Shift_7 (  ),
      .Dbg_Update_7 (  ),
      .Dbg_Rst_7 (  ),
      .Dbg_Clk_8 (  ),
      .Dbg_TDI_8 (  ),
      .Dbg_TDO_8 ( net_gnd0 ),
      .Dbg_Reg_En_8 (  ),
      .Dbg_Capture_8 (  ),
      .Dbg_Shift_8 (  ),
      .Dbg_Update_8 (  ),
      .Dbg_Rst_8 (  ),
      .Dbg_Clk_9 (  ),
      .Dbg_TDI_9 (  ),
      .Dbg_TDO_9 ( net_gnd0 ),
      .Dbg_Reg_En_9 (  ),
      .Dbg_Capture_9 (  ),
      .Dbg_Shift_9 (  ),
      .Dbg_Update_9 (  ),
      .Dbg_Rst_9 (  ),
      .Dbg_Clk_10 (  ),
      .Dbg_TDI_10 (  ),
      .Dbg_TDO_10 ( net_gnd0 ),
      .Dbg_Reg_En_10 (  ),
      .Dbg_Capture_10 (  ),
      .Dbg_Shift_10 (  ),
      .Dbg_Update_10 (  ),
      .Dbg_Rst_10 (  ),
      .Dbg_Clk_11 (  ),
      .Dbg_TDI_11 (  ),
      .Dbg_TDO_11 ( net_gnd0 ),
      .Dbg_Reg_En_11 (  ),
      .Dbg_Capture_11 (  ),
      .Dbg_Shift_11 (  ),
      .Dbg_Update_11 (  ),
      .Dbg_Rst_11 (  ),
      .Dbg_Clk_12 (  ),
      .Dbg_TDI_12 (  ),
      .Dbg_TDO_12 ( net_gnd0 ),
      .Dbg_Reg_En_12 (  ),
      .Dbg_Capture_12 (  ),
      .Dbg_Shift_12 (  ),
      .Dbg_Update_12 (  ),
      .Dbg_Rst_12 (  ),
      .Dbg_Clk_13 (  ),
      .Dbg_TDI_13 (  ),
      .Dbg_TDO_13 ( net_gnd0 ),
      .Dbg_Reg_En_13 (  ),
      .Dbg_Capture_13 (  ),
      .Dbg_Shift_13 (  ),
      .Dbg_Update_13 (  ),
      .Dbg_Rst_13 (  ),
      .Dbg_Clk_14 (  ),
      .Dbg_TDI_14 (  ),
      .Dbg_TDO_14 ( net_gnd0 ),
      .Dbg_Reg_En_14 (  ),
      .Dbg_Capture_14 (  ),
      .Dbg_Shift_14 (  ),
      .Dbg_Update_14 (  ),
      .Dbg_Rst_14 (  ),
      .Dbg_Clk_15 (  ),
      .Dbg_TDI_15 (  ),
      .Dbg_TDO_15 ( net_gnd0 ),
      .Dbg_Reg_En_15 (  ),
      .Dbg_Capture_15 (  ),
      .Dbg_Shift_15 (  ),
      .Dbg_Update_15 (  ),
      .Dbg_Rst_15 (  ),
      .Dbg_Clk_16 (  ),
      .Dbg_TDI_16 (  ),
      .Dbg_TDO_16 ( net_gnd0 ),
      .Dbg_Reg_En_16 (  ),
      .Dbg_Capture_16 (  ),
      .Dbg_Shift_16 (  ),
      .Dbg_Update_16 (  ),
      .Dbg_Rst_16 (  ),
      .Dbg_Clk_17 (  ),
      .Dbg_TDI_17 (  ),
      .Dbg_TDO_17 ( net_gnd0 ),
      .Dbg_Reg_En_17 (  ),
      .Dbg_Capture_17 (  ),
      .Dbg_Shift_17 (  ),
      .Dbg_Update_17 (  ),
      .Dbg_Rst_17 (  ),
      .Dbg_Clk_18 (  ),
      .Dbg_TDI_18 (  ),
      .Dbg_TDO_18 ( net_gnd0 ),
      .Dbg_Reg_En_18 (  ),
      .Dbg_Capture_18 (  ),
      .Dbg_Shift_18 (  ),
      .Dbg_Update_18 (  ),
      .Dbg_Rst_18 (  ),
      .Dbg_Clk_19 (  ),
      .Dbg_TDI_19 (  ),
      .Dbg_TDO_19 ( net_gnd0 ),
      .Dbg_Reg_En_19 (  ),
      .Dbg_Capture_19 (  ),
      .Dbg_Shift_19 (  ),
      .Dbg_Update_19 (  ),
      .Dbg_Rst_19 (  ),
      .Dbg_Clk_20 (  ),
      .Dbg_TDI_20 (  ),
      .Dbg_TDO_20 ( net_gnd0 ),
      .Dbg_Reg_En_20 (  ),
      .Dbg_Capture_20 (  ),
      .Dbg_Shift_20 (  ),
      .Dbg_Update_20 (  ),
      .Dbg_Rst_20 (  ),
      .Dbg_Clk_21 (  ),
      .Dbg_TDI_21 (  ),
      .Dbg_TDO_21 ( net_gnd0 ),
      .Dbg_Reg_En_21 (  ),
      .Dbg_Capture_21 (  ),
      .Dbg_Shift_21 (  ),
      .Dbg_Update_21 (  ),
      .Dbg_Rst_21 (  ),
      .Dbg_Clk_22 (  ),
      .Dbg_TDI_22 (  ),
      .Dbg_TDO_22 ( net_gnd0 ),
      .Dbg_Reg_En_22 (  ),
      .Dbg_Capture_22 (  ),
      .Dbg_Shift_22 (  ),
      .Dbg_Update_22 (  ),
      .Dbg_Rst_22 (  ),
      .Dbg_Clk_23 (  ),
      .Dbg_TDI_23 (  ),
      .Dbg_TDO_23 ( net_gnd0 ),
      .Dbg_Reg_En_23 (  ),
      .Dbg_Capture_23 (  ),
      .Dbg_Shift_23 (  ),
      .Dbg_Update_23 (  ),
      .Dbg_Rst_23 (  ),
      .Dbg_Clk_24 (  ),
      .Dbg_TDI_24 (  ),
      .Dbg_TDO_24 ( net_gnd0 ),
      .Dbg_Reg_En_24 (  ),
      .Dbg_Capture_24 (  ),
      .Dbg_Shift_24 (  ),
      .Dbg_Update_24 (  ),
      .Dbg_Rst_24 (  ),
      .Dbg_Clk_25 (  ),
      .Dbg_TDI_25 (  ),
      .Dbg_TDO_25 ( net_gnd0 ),
      .Dbg_Reg_En_25 (  ),
      .Dbg_Capture_25 (  ),
      .Dbg_Shift_25 (  ),
      .Dbg_Update_25 (  ),
      .Dbg_Rst_25 (  ),
      .Dbg_Clk_26 (  ),
      .Dbg_TDI_26 (  ),
      .Dbg_TDO_26 ( net_gnd0 ),
      .Dbg_Reg_En_26 (  ),
      .Dbg_Capture_26 (  ),
      .Dbg_Shift_26 (  ),
      .Dbg_Update_26 (  ),
      .Dbg_Rst_26 (  ),
      .Dbg_Clk_27 (  ),
      .Dbg_TDI_27 (  ),
      .Dbg_TDO_27 ( net_gnd0 ),
      .Dbg_Reg_En_27 (  ),
      .Dbg_Capture_27 (  ),
      .Dbg_Shift_27 (  ),
      .Dbg_Update_27 (  ),
      .Dbg_Rst_27 (  ),
      .Dbg_Clk_28 (  ),
      .Dbg_TDI_28 (  ),
      .Dbg_TDO_28 ( net_gnd0 ),
      .Dbg_Reg_En_28 (  ),
      .Dbg_Capture_28 (  ),
      .Dbg_Shift_28 (  ),
      .Dbg_Update_28 (  ),
      .Dbg_Rst_28 (  ),
      .Dbg_Clk_29 (  ),
      .Dbg_TDI_29 (  ),
      .Dbg_TDO_29 ( net_gnd0 ),
      .Dbg_Reg_En_29 (  ),
      .Dbg_Capture_29 (  ),
      .Dbg_Shift_29 (  ),
      .Dbg_Update_29 (  ),
      .Dbg_Rst_29 (  ),
      .Dbg_Clk_30 (  ),
      .Dbg_TDI_30 (  ),
      .Dbg_TDO_30 ( net_gnd0 ),
      .Dbg_Reg_En_30 (  ),
      .Dbg_Capture_30 (  ),
      .Dbg_Shift_30 (  ),
      .Dbg_Update_30 (  ),
      .Dbg_Rst_30 (  ),
      .Dbg_Clk_31 (  ),
      .Dbg_TDI_31 (  ),
      .Dbg_TDO_31 ( net_gnd0 ),
      .Dbg_Reg_En_31 (  ),
      .Dbg_Capture_31 (  ),
      .Dbg_Shift_31 (  ),
      .Dbg_Update_31 (  ),
      .Dbg_Rst_31 (  ),
      .bscan_tdi (  ),
      .bscan_reset (  ),
      .bscan_shift (  ),
      .bscan_update (  ),
      .bscan_capture (  ),
      .bscan_sel1 (  ),
      .bscan_drck1 (  ),
      .bscan_tdo1 ( net_gnd0 ),
      .bscan_ext_tdi ( net_gnd0 ),
      .bscan_ext_reset ( net_gnd0 ),
      .bscan_ext_shift ( net_gnd0 ),
      .bscan_ext_update ( net_gnd0 ),
      .bscan_ext_capture ( net_gnd0 ),
      .bscan_ext_sel ( net_gnd0 ),
      .bscan_ext_drck ( net_gnd0 ),
      .bscan_ext_tdo (  ),
      .Ext_JTAG_DRCK (  ),
      .Ext_JTAG_RESET (  ),
      .Ext_JTAG_SEL (  ),
      .Ext_JTAG_CAPTURE (  ),
      .Ext_JTAG_SHIFT (  ),
      .Ext_JTAG_UPDATE (  ),
      .Ext_JTAG_TDI (  ),
      .Ext_JTAG_TDO ( net_gnd0 )
    );

  microblaze_proc_sys_reset_0_wrapper
    proc_sys_reset_0 (
      .Slowest_sync_clk ( clk_50_0000MHz ),
      .Ext_Reset_In ( sys_rst_s ),
      .Aux_Reset_In ( net_gnd0 ),
      .MB_Debug_Sys_Rst ( Debug_SYS_Rst ),
      .Core_Reset_Req_0 ( net_gnd0 ),
      .Chip_Reset_Req_0 ( net_gnd0 ),
      .System_Reset_Req_0 ( net_gnd0 ),
      .Core_Reset_Req_1 ( net_gnd0 ),
      .Chip_Reset_Req_1 ( net_gnd0 ),
      .System_Reset_Req_1 ( net_gnd0 ),
      .Dcm_locked ( Dcm_all_locked ),
      .RstcPPCresetcore_0 (  ),
      .RstcPPCresetchip_0 (  ),
      .RstcPPCresetsys_0 (  ),
      .RstcPPCresetcore_1 (  ),
      .RstcPPCresetchip_1 (  ),
      .RstcPPCresetsys_1 (  ),
      .MB_Reset ( mb_reset ),
      .Bus_Struct_Reset ( sys_bus_reset[0:0] ),
      .Peripheral_Reset (  ),
      .Interconnect_aresetn (  ),
      .Peripheral_aresetn (  )
    );

  microblaze_xps_intc_0_wrapper
    xps_intc_0 (
      .SPLB_Clk ( clk_50_0000MHz ),
      .SPLB_Rst ( mb_plb_SPLB_Rst[2] ),
      .PLB_ABus ( mb_plb_PLB_ABus ),
      .PLB_PAValid ( mb_plb_PLB_PAValid ),
      .PLB_masterID ( mb_plb_PLB_masterID[0:0] ),
      .PLB_RNW ( mb_plb_PLB_RNW ),
      .PLB_BE ( mb_plb_PLB_BE ),
      .PLB_size ( mb_plb_PLB_size ),
      .PLB_type ( mb_plb_PLB_type ),
      .PLB_wrDBus ( mb_plb_PLB_wrDBus ),
      .PLB_UABus ( mb_plb_PLB_UABus ),
      .PLB_SAValid ( mb_plb_PLB_SAValid ),
      .PLB_rdPrim ( mb_plb_PLB_rdPrim[2] ),
      .PLB_wrPrim ( mb_plb_PLB_wrPrim[2] ),
      .PLB_abort ( mb_plb_PLB_abort ),
      .PLB_busLock ( mb_plb_PLB_busLock ),
      .PLB_MSize ( mb_plb_PLB_MSize ),
      .PLB_lockErr ( mb_plb_PLB_lockErr ),
      .PLB_wrBurst ( mb_plb_PLB_wrBurst ),
      .PLB_rdBurst ( mb_plb_PLB_rdBurst ),
      .PLB_wrPendReq ( mb_plb_PLB_wrPendReq ),
      .PLB_rdPendReq ( mb_plb_PLB_rdPendReq ),
      .PLB_wrPendPri ( mb_plb_PLB_wrPendPri ),
      .PLB_rdPendPri ( mb_plb_PLB_rdPendPri ),
      .PLB_reqPri ( mb_plb_PLB_reqPri ),
      .PLB_TAttribute ( mb_plb_PLB_TAttribute ),
      .Sl_addrAck ( mb_plb_Sl_addrAck[2] ),
      .Sl_SSize ( mb_plb_Sl_SSize[4:5] ),
      .Sl_wait ( mb_plb_Sl_wait[2] ),
      .Sl_rearbitrate ( mb_plb_Sl_rearbitrate[2] ),
      .Sl_wrDAck ( mb_plb_Sl_wrDAck[2] ),
      .Sl_wrComp ( mb_plb_Sl_wrComp[2] ),
      .Sl_rdDBus ( mb_plb_Sl_rdDBus[64:95] ),
      .Sl_rdDAck ( mb_plb_Sl_rdDAck[2] ),
      .Sl_rdComp ( mb_plb_Sl_rdComp[2] ),
      .Sl_MBusy ( mb_plb_Sl_MBusy[4:5] ),
      .Sl_MWrErr ( mb_plb_Sl_MWrErr[4:5] ),
      .Sl_MRdErr ( mb_plb_Sl_MRdErr[4:5] ),
      .Sl_wrBTerm ( mb_plb_Sl_wrBTerm[2] ),
      .Sl_rdWdAddr ( mb_plb_Sl_rdWdAddr[8:11] ),
      .Sl_rdBTerm ( mb_plb_Sl_rdBTerm[2] ),
      .Sl_MIRQ ( mb_plb_Sl_MIRQ[4:5] ),
      .Intr ( RS232_Interrupt[0:0] ),
      .Irq ( microblaze_0_Interrupt )
    );

  microblaze_plb_dac_0_wrapper
    plb_dac_0 (
      .SPLB_Clk ( clk_50_0000MHz ),
      .SPLB_Rst ( mb_plb_SPLB_Rst[3] ),
      .PLB_ABus ( mb_plb_PLB_ABus ),
      .PLB_UABus ( mb_plb_PLB_UABus ),
      .PLB_PAValid ( mb_plb_PLB_PAValid ),
      .PLB_SAValid ( mb_plb_PLB_SAValid ),
      .PLB_rdPrim ( mb_plb_PLB_rdPrim[3] ),
      .PLB_wrPrim ( mb_plb_PLB_wrPrim[3] ),
      .PLB_masterID ( mb_plb_PLB_masterID[0:0] ),
      .PLB_abort ( mb_plb_PLB_abort ),
      .PLB_busLock ( mb_plb_PLB_busLock ),
      .PLB_RNW ( mb_plb_PLB_RNW ),
      .PLB_BE ( mb_plb_PLB_BE ),
      .PLB_MSize ( mb_plb_PLB_MSize ),
      .PLB_size ( mb_plb_PLB_size ),
      .PLB_type ( mb_plb_PLB_type ),
      .PLB_lockErr ( mb_plb_PLB_lockErr ),
      .PLB_wrDBus ( mb_plb_PLB_wrDBus ),
      .PLB_wrBurst ( mb_plb_PLB_wrBurst ),
      .PLB_rdBurst ( mb_plb_PLB_rdBurst ),
      .PLB_wrPendReq ( mb_plb_PLB_wrPendReq ),
      .PLB_rdPendReq ( mb_plb_PLB_rdPendReq ),
      .PLB_wrPendPri ( mb_plb_PLB_wrPendPri ),
      .PLB_rdPendPri ( mb_plb_PLB_rdPendPri ),
      .PLB_reqPri ( mb_plb_PLB_reqPri ),
      .PLB_TAttribute ( mb_plb_PLB_TAttribute ),
      .Sl_addrAck ( mb_plb_Sl_addrAck[3] ),
      .Sl_SSize ( mb_plb_Sl_SSize[6:7] ),
      .Sl_wait ( mb_plb_Sl_wait[3] ),
      .Sl_rearbitrate ( mb_plb_Sl_rearbitrate[3] ),
      .Sl_wrDAck ( mb_plb_Sl_wrDAck[3] ),
      .Sl_wrComp ( mb_plb_Sl_wrComp[3] ),
      .Sl_wrBTerm ( mb_plb_Sl_wrBTerm[3] ),
      .Sl_rdDBus ( mb_plb_Sl_rdDBus[96:127] ),
      .Sl_rdWdAddr ( mb_plb_Sl_rdWdAddr[12:15] ),
      .Sl_rdDAck ( mb_plb_Sl_rdDAck[3] ),
      .Sl_rdComp ( mb_plb_Sl_rdComp[3] ),
      .Sl_rdBTerm ( mb_plb_Sl_rdBTerm[3] ),
      .Sl_MBusy ( mb_plb_Sl_MBusy[6:7] ),
      .Sl_MWrErr ( mb_plb_Sl_MWrErr[6:7] ),
      .Sl_MRdErr ( mb_plb_Sl_MRdErr[6:7] ),
      .Sl_MIRQ ( mb_plb_Sl_MIRQ[6:7] ),
      .S_Data ( plb_dac_0_S_Data ),
      .S_DCLKIO ( plb_dac_0_S_DCLKIO ),
      .S_Clkout ( plb_dac_0_S_Clkout ),
      .S_PinMD ( plb_dac_0_S_PinMD ),
      .S_ClkMD ( plb_dac_0_S_ClkMD ),
      .S_Format ( plb_dac_0_S_Format ),
      .S_PWRDN ( plb_dac_0_S_PWRDN )
    );

endmodule

