** Profile: "Plan A with Capacitors-Test High Freq"  [ F:\Programs\Verilog\FPGA_Group\test_br0101\analog\br0101_ad9715\br0101_ad9715-pspicefiles\plan a with capacitors\test high freq.sim ] 

** Creating circuit file "Test High Freq.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "F:/Academic/FPGA/BR0101/Development/DAC/model/ada4899.lib" 
* From [PSPICE NETLIST] section of G:\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.0.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 30us 10us 10ns 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Plan A with Capacitors.net" 


.END
